`timescale 1ns/ 1ps

module dsconv_block_batch_normalization_weights_memory(
    input  wire                clk,
    input  wire                rst,
    input  wire                start,
    input  wire        [2: 0]  layer_sel,  // 8
    input  wire        [3: 0]  filter_sel, // 16
    output reg  signed [17: 0] p,
    output reg  signed [35: 0] q,
    output reg                 ready
);
    reg signed [17: 0] ps [0: 7][0: 15];
    reg signed [35: 0] qs [0: 7][0: 15];

    initial begin
        ps[0][0]<=236; ps[0][1]<=172; ps[0][2]<=132; ps[0][3]<=166; ps[0][4]<=168; ps[0][5]<=154; ps[0][6]<=132; ps[0][7]<=249; ps[0][8]<=139; ps[0][9]<=425; ps[0][10]<=152; ps[0][11]<= 89; ps[0][12]<=236; ps[0][13]<=163; ps[0][14]<=198; ps[0][15]<=579; 
        ps[1][0]<=191; ps[1][1]<=186; ps[1][2]<=234; ps[1][3]<=150; ps[1][4]<=136; ps[1][5]<=123; ps[1][6]<=185; ps[1][7]<=133; ps[1][8]<=140; ps[1][9]<=191; ps[1][10]<=209; ps[1][11]<=175; ps[1][12]<=106; ps[1][13]<=231; ps[1][14]<=203; ps[1][15]<=200; 
        ps[2][0]<=246; ps[2][1]<=140; ps[2][2]<=172; ps[2][3]<=213; ps[2][4]<=230; ps[2][5]<=140; ps[2][6]<=201; ps[2][7]<=215; ps[2][8]<=144; ps[2][9]<=225; ps[2][10]<=154; ps[2][11]<=137; ps[2][12]<=486; ps[2][13]<=184; ps[2][14]<=106; ps[2][15]<=219; 
        ps[3][0]<=225; ps[3][1]<= 92; ps[3][2]<=490; ps[3][3]<=132; ps[3][4]<=318; ps[3][5]<=138; ps[3][6]<=303; ps[3][7]<=153; ps[3][8]<=226; ps[3][9]<=209; ps[3][10]<=199; ps[3][11]<=257; ps[3][12]<=168; ps[3][13]<=188; ps[3][14]<=261; ps[3][15]<=221; 
        ps[4][0]<=326; ps[4][1]<=241; ps[4][2]<=263; ps[4][3]<=330; ps[4][4]<=121; ps[4][5]<=351; ps[4][6]<=274; ps[4][7]<=361; ps[4][8]<=419; ps[4][9]<=280; ps[4][10]<=336; ps[4][11]<=164; ps[4][12]<=513; ps[4][13]<=173; ps[4][14]<=370; ps[4][15]<=517; 
        ps[5][0]<=208; ps[5][1]<=265; ps[5][2]<=222; ps[5][3]<=431; ps[5][4]<=180; ps[5][5]<=200; ps[5][6]<=425; ps[5][7]<=581; ps[5][8]<=217; ps[5][9]<=376; ps[5][10]<=295; ps[5][11]<=295; ps[5][12]<=107; ps[5][13]<=267; ps[5][14]<=501; ps[5][15]<=490; 
        ps[6][0]<=437; ps[6][1]<=146; ps[6][2]<=589; ps[6][3]<=524; ps[6][4]<=207; ps[6][5]<=453; ps[6][6]<=230; ps[6][7]<=208; ps[6][8]<=707; ps[6][9]<=375; ps[6][10]<=187; ps[6][11]<=173; ps[6][12]<=268; ps[6][13]<=293; ps[6][14]<=196; ps[6][15]<=143; 
        ps[7][0]<=119; ps[7][1]<= 57; ps[7][2]<= 43; ps[7][3]<= 81; ps[7][4]<= 77; ps[7][5]<= 79; ps[7][6]<= 65; ps[7][7]<= 79; ps[7][8]<= 95; ps[7][9]<= 54; ps[7][10]<=  0; ps[7][11]<= 74; ps[7][12]<= 53; ps[7][13]<=217; ps[7][14]<=173; ps[7][15]<= 67; 

        qs[0][0]<=-239327; qs[0][1]<=  12063; qs[0][2]<= -66655; qs[0][3]<=-186421; qs[0][4]<=-146331; qs[0][5]<=-163164; qs[0][6]<=-317053; qs[0][7]<=-213904; qs[0][8]<=-184505; qs[0][9]<=-221590; qs[0][10]<=-266562; qs[0][11]<=-147593; qs[0][12]<=-216496; qs[0][13]<=-209626; qs[0][14]<=-111305; qs[0][15]<=-432765; 
        qs[1][0]<=-182337; qs[1][1]<= -65071; qs[1][2]<=-239225; qs[1][3]<=-206252; qs[1][4]<=-183568; qs[1][5]<= -63007; qs[1][6]<= -69806; qs[1][7]<=-198324; qs[1][8]<= -94005; qs[1][9]<=-181681; qs[1][10]<=-183772; qs[1][11]<= -56093; qs[1][12]<= -68937; qs[1][13]<= -92047; qs[1][14]<=-269687; qs[1][15]<= -95759; 
        qs[2][0]<=-215624; qs[2][1]<=-157730; qs[2][2]<=-257839; qs[2][3]<= -72342; qs[2][4]<=-236647; qs[2][5]<= -95130; qs[2][6]<=-131875; qs[2][7]<=-243119; qs[2][8]<= -40168; qs[2][9]<=-239535; qs[2][10]<= -63345; qs[2][11]<=-186700; qs[2][12]<=-377536; qs[2][13]<=-205504; qs[2][14]<= -97008; qs[2][15]<=-356652; 
        qs[3][0]<=-213443; qs[3][1]<=    298; qs[3][2]<=-327019; qs[3][3]<=-107705; qs[3][4]<=-284009; qs[3][5]<= -18785; qs[3][6]<= -25144; qs[3][7]<=   9383; qs[3][8]<=-181302; qs[3][9]<=-286034; qs[3][10]<=-211413; qs[3][11]<= -26412; qs[3][12]<=-109279; qs[3][13]<=-364773; qs[3][14]<= -88984; qs[3][15]<=-211453; 
        qs[4][0]<=-146242; qs[4][1]<= -62590; qs[4][2]<=-161167; qs[4][3]<= -34877; qs[4][4]<=-125945; qs[4][5]<=-122515; qs[4][6]<= -52428; qs[4][7]<=-138221; qs[4][8]<= -79814; qs[4][9]<= -60503; qs[4][10]<=-141419; qs[4][11]<= -22962; qs[4][12]<=-197080; qs[4][13]<= -49508; qs[4][14]<=  -4018; qs[4][15]<=-110207; 
        qs[5][0]<=-236362; qs[5][1]<= -70321; qs[5][2]<=  -4949; qs[5][3]<= 110203; qs[5][4]<= -98666; qs[5][5]<=-125909; qs[5][6]<=-301350; qs[5][7]<=-163247; qs[5][8]<=  23081; qs[5][9]<=-115583; qs[5][10]<= -16336; qs[5][11]<=   8556; qs[5][12]<= -62175; qs[5][13]<=-101690; qs[5][14]<=-130276; qs[5][15]<=-125453; 
        qs[6][0]<=-140872; qs[6][1]<=  27677; qs[6][2]<=  74058; qs[6][3]<=-226021; qs[6][4]<= -35340; qs[6][5]<=-153929; qs[6][6]<=-108476; qs[6][7]<= -51247; qs[6][8]<= -32735; qs[6][9]<=  10768; qs[6][10]<= -46070; qs[6][11]<=-215627; qs[6][12]<=-121544; qs[6][13]<=-143107; qs[6][14]<= -12266; qs[6][15]<=  -6510; 
        qs[7][0]<=-178482; qs[7][1]<=-144889; qs[7][2]<= -21921; qs[7][3]<=-222833; qs[7][4]<=-246133; qs[7][5]<=-193177; qs[7][6]<=-140128; qs[7][7]<= -90629; qs[7][8]<= -69026; qs[7][9]<=-217123; qs[7][10]<=    471; qs[7][11]<=-218205; qs[7][12]<=-152177; qs[7][13]<=-112706; qs[7][14]<=-155701; qs[7][15]<=-188089; 
    end

    always@(posedge clk) begin
        if(rst) begin
            p    <=0;
            q    <=0;
            ready<=0;
        end else if(start) begin
            p    <=ps[layer_sel][filter_sel];
            q    <=qs[layer_sel][filter_sel];
            ready<=1;
        end
    end
endmodule