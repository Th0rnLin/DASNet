`timescale 1ns/ 1ps

module dsconv_block_depthwise_weights_memory(
    input  wire                clk,
    input  wire                rst,
    input  wire                start,
    input  wire        [2: 0]  layer_sel,  // 8
    input  wire        [3: 0]  filter_sel, // 16
    output reg  signed [17: 0] w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48,
    output reg                 ready
);
    reg signed [17: 0] ws [7: 0][0: 15][0: 48];

    initial begin
        ws[0][0 ][0]<=  28; ws[0][0 ][1]<=  39; ws[0][0 ][2]<=-147; ws[0][0 ][3]<= -85; ws[0][0 ][4]<=  27; ws[0][0 ][5]<= 101; ws[0][0 ][6]<=  99; ws[0][0 ][7]<=  44; ws[0][0 ][8]<=  88; ws[0][0 ][9]<= -50; ws[0][0 ][10]<= -35; ws[0][0 ][11]<=  98; ws[0][0 ][12]<= 230; ws[0][0 ][13]<=  41; ws[0][0 ][14]<=  28; ws[0][0 ][15]<= -14; ws[0][0 ][16]<=  -7; ws[0][0 ][17]<=  30; ws[0][0 ][18]<= 173; ws[0][0 ][19]<= 238; ws[0][0 ][20]<=  17; ws[0][0 ][21]<= -20; ws[0][0 ][22]<=  60; ws[0][0 ][23]<=  39; ws[0][0 ][24]<=   0; ws[0][0 ][25]<= 100; ws[0][0 ][26]<= 156; ws[0][0 ][27]<= -43; ws[0][0 ][28]<=  50; ws[0][0 ][29]<=  14; ws[0][0 ][30]<= -28; ws[0][0 ][31]<= -20; ws[0][0 ][32]<= -42; ws[0][0 ][33]<=  41; ws[0][0 ][34]<= -49; ws[0][0 ][35]<=  45; ws[0][0 ][36]<=  24; ws[0][0 ][37]<= -36; ws[0][0 ][38]<= -74; ws[0][0 ][39]<=-104; ws[0][0 ][40]<= -25; ws[0][0 ][41]<= -66; ws[0][0 ][42]<=  26; ws[0][0 ][43]<=-123; ws[0][0 ][44]<=-211; ws[0][0 ][45]<=-232; ws[0][0 ][46]<=-253; ws[0][0 ][47]<=-165; ws[0][0 ][48]<=-117;
        ws[0][1 ][0]<=  23; ws[0][1 ][1]<=  10; ws[0][1 ][2]<=  39; ws[0][1 ][3]<=  23; ws[0][1 ][4]<=  54; ws[0][1 ][5]<=  34; ws[0][1 ][6]<=  16; ws[0][1 ][7]<=  34; ws[0][1 ][8]<=  34; ws[0][1 ][9]<=  17; ws[0][1 ][10]<=  95; ws[0][1 ][11]<= 102; ws[0][1 ][12]<=  95; ws[0][1 ][13]<=  98; ws[0][1 ][14]<=  50; ws[0][1 ][15]<=  60; ws[0][1 ][16]<=  67; ws[0][1 ][17]<=  19; ws[0][1 ][18]<=  86; ws[0][1 ][19]<=  58; ws[0][1 ][20]<=  51; ws[0][1 ][21]<=  -3; ws[0][1 ][22]<=  81; ws[0][1 ][23]<=  33; ws[0][1 ][24]<=  76; ws[0][1 ][25]<=  56; ws[0][1 ][26]<=  18; ws[0][1 ][27]<=  44; ws[0][1 ][28]<=   6; ws[0][1 ][29]<=  57; ws[0][1 ][30]<=  97; ws[0][1 ][31]<=  97; ws[0][1 ][32]<=  27; ws[0][1 ][33]<=  81; ws[0][1 ][34]<=  75; ws[0][1 ][35]<=  -9; ws[0][1 ][36]<=  20; ws[0][1 ][37]<=  40; ws[0][1 ][38]<=  66; ws[0][1 ][39]<=  71; ws[0][1 ][40]<=  32; ws[0][1 ][41]<=  85; ws[0][1 ][42]<=  61; ws[0][1 ][43]<= -20; ws[0][1 ][44]<=  59; ws[0][1 ][45]<=  25; ws[0][1 ][46]<=  50; ws[0][1 ][47]<=  68; ws[0][1 ][48]<=  50;
        ws[0][2 ][0]<=   4; ws[0][2 ][1]<=  99; ws[0][2 ][2]<= -44; ws[0][2 ][3]<=-142; ws[0][2 ][4]<= -79; ws[0][2 ][5]<=  -8; ws[0][2 ][6]<= -55; ws[0][2 ][7]<=  81; ws[0][2 ][8]<=  81; ws[0][2 ][9]<=-119; ws[0][2 ][10]<=-214; ws[0][2 ][11]<=-129; ws[0][2 ][12]<= -36; ws[0][2 ][13]<= -39; ws[0][2 ][14]<= 141; ws[0][2 ][15]<= 152; ws[0][2 ][16]<= -75; ws[0][2 ][17]<=-199; ws[0][2 ][18]<=-139; ws[0][2 ][19]<= -40; ws[0][2 ][20]<= -76; ws[0][2 ][21]<= 194; ws[0][2 ][22]<= 181; ws[0][2 ][23]<= -82; ws[0][2 ][24]<=-138; ws[0][2 ][25]<= -15; ws[0][2 ][26]<=  99; ws[0][2 ][27]<= -85; ws[0][2 ][28]<= 130; ws[0][2 ][29]<=  78; ws[0][2 ][30]<=  34; ws[0][2 ][31]<=-101; ws[0][2 ][32]<=  -9; ws[0][2 ][33]<= 102; ws[0][2 ][34]<=-128; ws[0][2 ][35]<=  36; ws[0][2 ][36]<= 111; ws[0][2 ][37]<= 150; ws[0][2 ][38]<=  15; ws[0][2 ][39]<=  83; ws[0][2 ][40]<=  59; ws[0][2 ][41]<= -75; ws[0][2 ][42]<=-135; ws[0][2 ][43]<=  78; ws[0][2 ][44]<= 142; ws[0][2 ][45]<=  85; ws[0][2 ][46]<=  30; ws[0][2 ][47]<=  -8; ws[0][2 ][48]<= -74;
        ws[0][3 ][0]<=-124; ws[0][3 ][1]<= -43; ws[0][3 ][2]<=  31; ws[0][3 ][3]<=  23; ws[0][3 ][4]<= -84; ws[0][3 ][5]<=-217; ws[0][3 ][6]<=-103; ws[0][3 ][7]<=-143; ws[0][3 ][8]<=-116; ws[0][3 ][9]<= -20; ws[0][3 ][10]<=  57; ws[0][3 ][11]<=-116; ws[0][3 ][12]<=-202; ws[0][3 ][13]<= -77; ws[0][3 ][14]<= -60; ws[0][3 ][15]<=-112; ws[0][3 ][16]<= -43; ws[0][3 ][17]<=  39; ws[0][3 ][18]<= -45; ws[0][3 ][19]<=-219; ws[0][3 ][20]<= -46; ws[0][3 ][21]<=  59; ws[0][3 ][22]<=-116; ws[0][3 ][23]<=  -1; ws[0][3 ][24]<=  74; ws[0][3 ][25]<= -34; ws[0][3 ][26]<=-154; ws[0][3 ][27]<= -40; ws[0][3 ][28]<= 118; ws[0][3 ][29]<=  -8; ws[0][3 ][30]<=  76; ws[0][3 ][31]<= 132; ws[0][3 ][32]<=  81; ws[0][3 ][33]<= -18; ws[0][3 ][34]<=  -1; ws[0][3 ][35]<=  26; ws[0][3 ][36]<= -41; ws[0][3 ][37]<=  67; ws[0][3 ][38]<= 164; ws[0][3 ][39]<= 158; ws[0][3 ][40]<= 128; ws[0][3 ][41]<=  73; ws[0][3 ][42]<= -47; ws[0][3 ][43]<=  29; ws[0][3 ][44]<= 122; ws[0][3 ][45]<= 221; ws[0][3 ][46]<= 200; ws[0][3 ][47]<= 171; ws[0][3 ][48]<= 164;
        ws[0][4 ][0]<= -57; ws[0][4 ][1]<= -41; ws[0][4 ][2]<= -87; ws[0][4 ][3]<= -40; ws[0][4 ][4]<= 196; ws[0][4 ][5]<= 227; ws[0][4 ][6]<= 278; ws[0][4 ][7]<= -59; ws[0][4 ][8]<=  17; ws[0][4 ][9]<= -92; ws[0][4 ][10]<= -27; ws[0][4 ][11]<=  88; ws[0][4 ][12]<= 182; ws[0][4 ][13]<= 152; ws[0][4 ][14]<=-117; ws[0][4 ][15]<=  -7; ws[0][4 ][16]<= -75; ws[0][4 ][17]<=-123; ws[0][4 ][18]<= -14; ws[0][4 ][19]<= 138; ws[0][4 ][20]<=  60; ws[0][4 ][21]<=-133; ws[0][4 ][22]<=  -5; ws[0][4 ][23]<= -55; ws[0][4 ][24]<=-117; ws[0][4 ][25]<= -81; ws[0][4 ][26]<=  69; ws[0][4 ][27]<=  18; ws[0][4 ][28]<=-154; ws[0][4 ][29]<= -20; ws[0][4 ][30]<= -21; ws[0][4 ][31]<=-119; ws[0][4 ][32]<=-109; ws[0][4 ][33]<= -34; ws[0][4 ][34]<= 100; ws[0][4 ][35]<=-141; ws[0][4 ][36]<=  -7; ws[0][4 ][37]<= -16; ws[0][4 ][38]<= -72; ws[0][4 ][39]<= -14; ws[0][4 ][40]<= 125; ws[0][4 ][41]<= 121; ws[0][4 ][42]<=-139; ws[0][4 ][43]<= -88; ws[0][4 ][44]<= -19; ws[0][4 ][45]<=  34; ws[0][4 ][46]<=  79; ws[0][4 ][47]<= 202; ws[0][4 ][48]<= 214;
        ws[0][5 ][0]<=  86; ws[0][5 ][1]<= -19; ws[0][5 ][2]<= -55; ws[0][5 ][3]<=  97; ws[0][5 ][4]<= 164; ws[0][5 ][5]<= 153; ws[0][5 ][6]<=  80; ws[0][5 ][7]<=  96; ws[0][5 ][8]<=-194; ws[0][5 ][9]<=-202; ws[0][5 ][10]<= -51; ws[0][5 ][11]<= 103; ws[0][5 ][12]<=  66; ws[0][5 ][13]<= -59; ws[0][5 ][14]<=  63; ws[0][5 ][15]<=-202; ws[0][5 ][16]<=-234; ws[0][5 ][17]<= -25; ws[0][5 ][18]<=  83; ws[0][5 ][19]<=  42; ws[0][5 ][20]<= -88; ws[0][5 ][21]<=  81; ws[0][5 ][22]<=-146; ws[0][5 ][23]<=-120; ws[0][5 ][24]<= -26; ws[0][5 ][25]<=  84; ws[0][5 ][26]<=  14; ws[0][5 ][27]<=-126; ws[0][5 ][28]<=  92; ws[0][5 ][29]<= -56; ws[0][5 ][30]<=-112; ws[0][5 ][31]<=  42; ws[0][5 ][32]<= 141; ws[0][5 ][33]<=  39; ws[0][5 ][34]<=-154; ws[0][5 ][35]<=  52; ws[0][5 ][36]<= -68; ws[0][5 ][37]<=-102; ws[0][5 ][38]<= -18; ws[0][5 ][39]<=  68; ws[0][5 ][40]<=  57; ws[0][5 ][41]<= -60; ws[0][5 ][42]<= 113; ws[0][5 ][43]<=  21; ws[0][5 ][44]<= -19; ws[0][5 ][45]<=  45; ws[0][5 ][46]<=  96; ws[0][5 ][47]<=  65; ws[0][5 ][48]<= -73;
        ws[0][6 ][0]<=  64; ws[0][6 ][1]<=  43; ws[0][6 ][2]<= 107; ws[0][6 ][3]<= 179; ws[0][6 ][4]<= 327; ws[0][6 ][5]<= 179; ws[0][6 ][6]<= 134; ws[0][6 ][7]<=  89; ws[0][6 ][8]<=  75; ws[0][6 ][9]<= 141; ws[0][6 ][10]<= 206; ws[0][6 ][11]<= 258; ws[0][6 ][12]<= 155; ws[0][6 ][13]<=  98; ws[0][6 ][14]<=  10; ws[0][6 ][15]<=  24; ws[0][6 ][16]<=  46; ws[0][6 ][17]<= 148; ws[0][6 ][18]<= 178; ws[0][6 ][19]<= 143; ws[0][6 ][20]<= 104; ws[0][6 ][21]<= -48; ws[0][6 ][22]<= -58; ws[0][6 ][23]<=  14; ws[0][6 ][24]<=  29; ws[0][6 ][25]<= 108; ws[0][6 ][26]<= 112; ws[0][6 ][27]<= 103; ws[0][6 ][28]<= -16; ws[0][6 ][29]<= -12; ws[0][6 ][30]<= -67; ws[0][6 ][31]<=  50; ws[0][6 ][32]<= 103; ws[0][6 ][33]<= 142; ws[0][6 ][34]<=  51; ws[0][6 ][35]<= -47; ws[0][6 ][36]<=   8; ws[0][6 ][37]<=   6; ws[0][6 ][38]<=  15; ws[0][6 ][39]<= 182; ws[0][6 ][40]<= 169; ws[0][6 ][41]<= 102; ws[0][6 ][42]<=  29; ws[0][6 ][43]<=  34; ws[0][6 ][44]<=  -9; ws[0][6 ][45]<= 147; ws[0][6 ][46]<= 242; ws[0][6 ][47]<= 205; ws[0][6 ][48]<= 121;
        ws[0][7 ][0]<=   3; ws[0][7 ][1]<=   1; ws[0][7 ][2]<= -40; ws[0][7 ][3]<= -28; ws[0][7 ][4]<=  59; ws[0][7 ][5]<=  81; ws[0][7 ][6]<= 141; ws[0][7 ][7]<=  -1; ws[0][7 ][8]<=  77; ws[0][7 ][9]<=  42; ws[0][7 ][10]<= -56; ws[0][7 ][11]<= -66; ws[0][7 ][12]<= -40; ws[0][7 ][13]<= -20; ws[0][7 ][14]<= -18; ws[0][7 ][15]<=  11; ws[0][7 ][16]<=  65; ws[0][7 ][17]<= -58; ws[0][7 ][18]<=-180; ws[0][7 ][19]<=-169; ws[0][7 ][20]<=-143; ws[0][7 ][21]<=  24; ws[0][7 ][22]<=  63; ws[0][7 ][23]<=  75; ws[0][7 ][24]<= -71; ws[0][7 ][25]<=-248; ws[0][7 ][26]<=-265; ws[0][7 ][27]<=-164; ws[0][7 ][28]<=  -6; ws[0][7 ][29]<=  26; ws[0][7 ][30]<=  34; ws[0][7 ][31]<= -41; ws[0][7 ][32]<=-250; ws[0][7 ][33]<=-179; ws[0][7 ][34]<= -95; ws[0][7 ][35]<=  65; ws[0][7 ][36]<=  31; ws[0][7 ][37]<=  38; ws[0][7 ][38]<=  -5; ws[0][7 ][39]<=-195; ws[0][7 ][40]<=-235; ws[0][7 ][41]<= -64; ws[0][7 ][42]<= -39; ws[0][7 ][43]<= -48; ws[0][7 ][44]<= -16; ws[0][7 ][45]<=  -3; ws[0][7 ][46]<=-207; ws[0][7 ][47]<=-270; ws[0][7 ][48]<=-136;
        ws[0][8 ][0]<= 137; ws[0][8 ][1]<=  31; ws[0][8 ][2]<= -27; ws[0][8 ][3]<=  89; ws[0][8 ][4]<= 150; ws[0][8 ][5]<=  93; ws[0][8 ][6]<= 228; ws[0][8 ][7]<= 132; ws[0][8 ][8]<=  68; ws[0][8 ][9]<=  56; ws[0][8 ][10]<=  65; ws[0][8 ][11]<=  86; ws[0][8 ][12]<=  84; ws[0][8 ][13]<= 167; ws[0][8 ][14]<=  45; ws[0][8 ][15]<= 109; ws[0][8 ][16]<=  47; ws[0][8 ][17]<=  11; ws[0][8 ][18]<=  50; ws[0][8 ][19]<=  66; ws[0][8 ][20]<= 111; ws[0][8 ][21]<=  66; ws[0][8 ][22]<=  93; ws[0][8 ][23]<=  52; ws[0][8 ][24]<=   3; ws[0][8 ][25]<= -26; ws[0][8 ][26]<=  65; ws[0][8 ][27]<=  65; ws[0][8 ][28]<=  56; ws[0][8 ][29]<=  58; ws[0][8 ][30]<=  99; ws[0][8 ][31]<=  24; ws[0][8 ][32]<= -38; ws[0][8 ][33]<=   7; ws[0][8 ][34]<= -11; ws[0][8 ][35]<=  48; ws[0][8 ][36]<=  38; ws[0][8 ][37]<= 172; ws[0][8 ][38]<=  78; ws[0][8 ][39]<=   8; ws[0][8 ][40]<=  44; ws[0][8 ][41]<=  62; ws[0][8 ][42]<= -69; ws[0][8 ][43]<=  30; ws[0][8 ][44]<= 177; ws[0][8 ][45]<= 138; ws[0][8 ][46]<=  77; ws[0][8 ][47]<=  33; ws[0][8 ][48]<=  80;
        ws[0][9 ][0]<= -23; ws[0][9 ][1]<=  97; ws[0][9 ][2]<=   1; ws[0][9 ][3]<= -93; ws[0][9 ][4]<=-128; ws[0][9 ][5]<=-195; ws[0][9 ][6]<=-102; ws[0][9 ][7]<=  14; ws[0][9 ][8]<= 120; ws[0][9 ][9]<=  43; ws[0][9 ][10]<=-124; ws[0][9 ][11]<= -72; ws[0][9 ][12]<= -80; ws[0][9 ][13]<= -45; ws[0][9 ][14]<= -89; ws[0][9 ][15]<= 125; ws[0][9 ][16]<= -48; ws[0][9 ][17]<=-101; ws[0][9 ][18]<=   1; ws[0][9 ][19]<= -62; ws[0][9 ][20]<= -81; ws[0][9 ][21]<=-115; ws[0][9 ][22]<= -29; ws[0][9 ][23]<=-139; ws[0][9 ][24]<=-235; ws[0][9 ][25]<=   6; ws[0][9 ][26]<=  54; ws[0][9 ][27]<=  14; ws[0][9 ][28]<= -59; ws[0][9 ][29]<= -56; ws[0][9 ][30]<=-133; ws[0][9 ][31]<=-225; ws[0][9 ][32]<= -60; ws[0][9 ][33]<=  -1; ws[0][9 ][34]<=  26; ws[0][9 ][35]<=  65; ws[0][9 ][36]<= 104; ws[0][9 ][37]<= -35; ws[0][9 ][38]<=-112; ws[0][9 ][39]<=  16; ws[0][9 ][40]<=  72; ws[0][9 ][41]<= 115; ws[0][9 ][42]<= 163; ws[0][9 ][43]<= 210; ws[0][9 ][44]<=  73; ws[0][9 ][45]<= -63; ws[0][9 ][46]<=  74; ws[0][9 ][47]<= 221; ws[0][9 ][48]<= 232;
        ws[0][10][0]<= -95; ws[0][10][1]<= -17; ws[0][10][2]<=-130; ws[0][10][3]<=-104; ws[0][10][4]<= -66; ws[0][10][5]<= -65; ws[0][10][6]<=  41; ws[0][10][7]<= -84; ws[0][10][8]<= -84; ws[0][10][9]<=-102; ws[0][10][10]<= -57; ws[0][10][11]<=  54; ws[0][10][12]<=  29; ws[0][10][13]<= -30; ws[0][10][14]<= -53; ws[0][10][15]<=-134; ws[0][10][16]<= -69; ws[0][10][17]<=   7; ws[0][10][18]<= 160; ws[0][10][19]<= 141; ws[0][10][20]<= -28; ws[0][10][21]<=  25; ws[0][10][22]<= -69; ws[0][10][23]<= -22; ws[0][10][24]<= 157; ws[0][10][25]<= 197; ws[0][10][26]<= 158; ws[0][10][27]<=-145; ws[0][10][28]<=  32; ws[0][10][29]<=  58; ws[0][10][30]<=  86; ws[0][10][31]<= 174; ws[0][10][32]<= 169; ws[0][10][33]<=  91; ws[0][10][34]<=-201; ws[0][10][35]<=  56; ws[0][10][36]<=  58; ws[0][10][37]<= 115; ws[0][10][38]<=  95; ws[0][10][39]<=  75; ws[0][10][40]<=  50; ws[0][10][41]<= -77; ws[0][10][42]<=-103; ws[0][10][43]<= -39; ws[0][10][44]<=  12; ws[0][10][45]<=  51; ws[0][10][46]<= -14; ws[0][10][47]<=   9; ws[0][10][48]<= -28;
        ws[0][11][0]<= -23; ws[0][11][1]<=  -8; ws[0][11][2]<=   7; ws[0][11][3]<=  37; ws[0][11][4]<= -34; ws[0][11][5]<=-107; ws[0][11][6]<= -25; ws[0][11][7]<= -70; ws[0][11][8]<=  -8; ws[0][11][9]<=  25; ws[0][11][10]<= -21; ws[0][11][11]<= -70; ws[0][11][12]<= -86; ws[0][11][13]<= -86; ws[0][11][14]<= -52; ws[0][11][15]<=   5; ws[0][11][16]<=  10; ws[0][11][17]<= -57; ws[0][11][18]<= -44; ws[0][11][19]<=-133; ws[0][11][20]<=-107; ws[0][11][21]<= -22; ws[0][11][22]<= -41; ws[0][11][23]<=  10; ws[0][11][24]<= -16; ws[0][11][25]<= -85; ws[0][11][26]<= -45; ws[0][11][27]<= -76; ws[0][11][28]<=-101; ws[0][11][29]<= -54; ws[0][11][30]<=   6; ws[0][11][31]<=  21; ws[0][11][32]<= -23; ws[0][11][33]<= -85; ws[0][11][34]<= -63; ws[0][11][35]<=-119; ws[0][11][36]<=  -1; ws[0][11][37]<= -18; ws[0][11][38]<=  15; ws[0][11][39]<= -34; ws[0][11][40]<= -50; ws[0][11][41]<= -42; ws[0][11][42]<=-115; ws[0][11][43]<= -58; ws[0][11][44]<=  42; ws[0][11][45]<= -16; ws[0][11][46]<=  18; ws[0][11][47]<= -48; ws[0][11][48]<=  46;
        ws[0][12][0]<= -73; ws[0][12][1]<=  40; ws[0][12][2]<=  44; ws[0][12][3]<= -61; ws[0][12][4]<= -26; ws[0][12][5]<=  39; ws[0][12][6]<=   5; ws[0][12][7]<= -15; ws[0][12][8]<= 134; ws[0][12][9]<=  96; ws[0][12][10]<= -81; ws[0][12][11]<=-122; ws[0][12][12]<=  -4; ws[0][12][13]<= -34; ws[0][12][14]<=  69; ws[0][12][15]<= 148; ws[0][12][16]<=  39; ws[0][12][17]<=-293; ws[0][12][18]<=-369; ws[0][12][19]<= -79; ws[0][12][20]<=-125; ws[0][12][21]<=  40; ws[0][12][22]<= 131; ws[0][12][23]<= -89; ws[0][12][24]<=-378; ws[0][12][25]<=-433; ws[0][12][26]<=-117; ws[0][12][27]<= -58; ws[0][12][28]<= -34; ws[0][12][29]<=  17; ws[0][12][30]<= -43; ws[0][12][31]<=-301; ws[0][12][32]<=-339; ws[0][12][33]<= -56; ws[0][12][34]<= -75; ws[0][12][35]<=  15; ws[0][12][36]<=  55; ws[0][12][37]<= -25; ws[0][12][38]<= -87; ws[0][12][39]<=-113; ws[0][12][40]<=  34; ws[0][12][41]<= -71; ws[0][12][42]<=  16; ws[0][12][43]<=  45; ws[0][12][44]<=  46; ws[0][12][45]<= -27; ws[0][12][46]<=  51; ws[0][12][47]<=  25; ws[0][12][48]<= -61;
        ws[0][13][0]<=  13; ws[0][13][1]<=-117; ws[0][13][2]<=-118; ws[0][13][3]<=-127; ws[0][13][4]<=  37; ws[0][13][5]<=  74; ws[0][13][6]<=  -9; ws[0][13][7]<= -10; ws[0][13][8]<= -41; ws[0][13][9]<= -86; ws[0][13][10]<= -75; ws[0][13][11]<= 103; ws[0][13][12]<= 154; ws[0][13][13]<=  92; ws[0][13][14]<=   8; ws[0][13][15]<=  19; ws[0][13][16]<= -27; ws[0][13][17]<=  -3; ws[0][13][18]<=  17; ws[0][13][19]<=  73; ws[0][13][20]<=  -8; ws[0][13][21]<= -48; ws[0][13][22]<=  83; ws[0][13][23]<=  26; ws[0][13][24]<= -56; ws[0][13][25]<= -38; ws[0][13][26]<=  71; ws[0][13][27]<=  40; ws[0][13][28]<= -40; ws[0][13][29]<=  44; ws[0][13][30]<=  57; ws[0][13][31]<= -30; ws[0][13][32]<= -23; ws[0][13][33]<= -25; ws[0][13][34]<= -76; ws[0][13][35]<=   7; ws[0][13][36]<=  49; ws[0][13][37]<= -44; ws[0][13][38]<= -87; ws[0][13][39]<= -60; ws[0][13][40]<=-129; ws[0][13][41]<=-136; ws[0][13][42]<= 135; ws[0][13][43]<= 107; ws[0][13][44]<= -67; ws[0][13][45]<=-140; ws[0][13][46]<= -97; ws[0][13][47]<=-174; ws[0][13][48]<=-198;
        ws[0][14][0]<=  53; ws[0][14][1]<=  78; ws[0][14][2]<=  22; ws[0][14][3]<= -25; ws[0][14][4]<=  23; ws[0][14][5]<=  38; ws[0][14][6]<=-146; ws[0][14][7]<=  94; ws[0][14][8]<=  33; ws[0][14][9]<= -14; ws[0][14][10]<=  -6; ws[0][14][11]<=  83; ws[0][14][12]<= 128; ws[0][14][13]<= -92; ws[0][14][14]<=  72; ws[0][14][15]<=  91; ws[0][14][16]<=  17; ws[0][14][17]<= -28; ws[0][14][18]<=  55; ws[0][14][19]<=  91; ws[0][14][20]<=   0; ws[0][14][21]<=  71; ws[0][14][22]<= 110; ws[0][14][23]<=  25; ws[0][14][24]<= -20; ws[0][14][25]<=  52; ws[0][14][26]<=  85; ws[0][14][27]<=  24; ws[0][14][28]<=  56; ws[0][14][29]<= 153; ws[0][14][30]<=  10; ws[0][14][31]<= -19; ws[0][14][32]<= -24; ws[0][14][33]<=  95; ws[0][14][34]<=  -6; ws[0][14][35]<=  81; ws[0][14][36]<= 170; ws[0][14][37]<=  63; ws[0][14][38]<= -22; ws[0][14][39]<=   0; ws[0][14][40]<=  63; ws[0][14][41]<= -37; ws[0][14][42]<= 110; ws[0][14][43]<= 138; ws[0][14][44]<=  67; ws[0][14][45]<=-105; ws[0][14][46]<= -80; ws[0][14][47]<= -24; ws[0][14][48]<= -74;
        ws[0][15][0]<= -30; ws[0][15][1]<=  38; ws[0][15][2]<=  39; ws[0][15][3]<=   6; ws[0][15][4]<=  81; ws[0][15][5]<=  86; ws[0][15][6]<=  72; ws[0][15][7]<=  29; ws[0][15][8]<=  43; ws[0][15][9]<=  63; ws[0][15][10]<= -26; ws[0][15][11]<=  30; ws[0][15][12]<=  88; ws[0][15][13]<=  40; ws[0][15][14]<=  37; ws[0][15][15]<=  65; ws[0][15][16]<=  55; ws[0][15][17]<=  10; ws[0][15][18]<=  10; ws[0][15][19]<=  -6; ws[0][15][20]<=  19; ws[0][15][21]<=  28; ws[0][15][22]<= 139; ws[0][15][23]<= 125; ws[0][15][24]<=  34; ws[0][15][25]<=   0; ws[0][15][26]<=  29; ws[0][15][27]<=  25; ws[0][15][28]<= -24; ws[0][15][29]<= 112; ws[0][15][30]<=  64; ws[0][15][31]<=  44; ws[0][15][32]<= -35; ws[0][15][33]<=  20; ws[0][15][34]<=  -5; ws[0][15][35]<= -23; ws[0][15][36]<= 117; ws[0][15][37]<= 114; ws[0][15][38]<=  57; ws[0][15][39]<= -34; ws[0][15][40]<=   0; ws[0][15][41]<=  -8; ws[0][15][42]<= -78; ws[0][15][43]<=  46; ws[0][15][44]<= 129; ws[0][15][45]<=  58; ws[0][15][46]<=  40; ws[0][15][47]<=  -1; ws[0][15][48]<=  41;

        ws[1][0 ][0]<=  75; ws[1][0 ][1]<= -28; ws[1][0 ][2]<=  38; ws[1][0 ][3]<=  64; ws[1][0 ][4]<= 120; ws[1][0 ][5]<= 144; ws[1][0 ][6]<=  46; ws[1][0 ][7]<=  63; ws[1][0 ][8]<=  35; ws[1][0 ][9]<=  -8; ws[1][0 ][10]<=  61; ws[1][0 ][11]<=  68; ws[1][0 ][12]<=  59; ws[1][0 ][13]<=  36; ws[1][0 ][14]<= 143; ws[1][0 ][15]<=  30; ws[1][0 ][16]<= -47; ws[1][0 ][17]<=  39; ws[1][0 ][18]<=  51; ws[1][0 ][19]<=  74; ws[1][0 ][20]<=  78; ws[1][0 ][21]<= 133; ws[1][0 ][22]<=  68; ws[1][0 ][23]<= -39; ws[1][0 ][24]<= -45; ws[1][0 ][25]<=  50; ws[1][0 ][26]<=  58; ws[1][0 ][27]<=  74; ws[1][0 ][28]<=  91; ws[1][0 ][29]<=  70; ws[1][0 ][30]<=  23; ws[1][0 ][31]<= -28; ws[1][0 ][32]<=  51; ws[1][0 ][33]<=  94; ws[1][0 ][34]<=  77; ws[1][0 ][35]<= 107; ws[1][0 ][36]<=  16; ws[1][0 ][37]<= -35; ws[1][0 ][38]<=   4; ws[1][0 ][39]<=  -7; ws[1][0 ][40]<=  96; ws[1][0 ][41]<=  93; ws[1][0 ][42]<=  38; ws[1][0 ][43]<=   6; ws[1][0 ][44]<= -88; ws[1][0 ][45]<= -13; ws[1][0 ][46]<= -16; ws[1][0 ][47]<=  31; ws[1][0 ][48]<=  63;
        ws[1][1 ][0]<=  54; ws[1][1 ][1]<=  -7; ws[1][1 ][2]<=  68; ws[1][1 ][3]<= 132; ws[1][1 ][4]<=  73; ws[1][1 ][5]<=  14; ws[1][1 ][6]<= -19; ws[1][1 ][7]<= -25; ws[1][1 ][8]<=  80; ws[1][1 ][9]<= 131; ws[1][1 ][10]<=  46; ws[1][1 ][11]<=  -2; ws[1][1 ][12]<= -57; ws[1][1 ][13]<= -84; ws[1][1 ][14]<= -93; ws[1][1 ][15]<= 138; ws[1][1 ][16]<=  90; ws[1][1 ][17]<= -29; ws[1][1 ][18]<=-168; ws[1][1 ][19]<=-143; ws[1][1 ][20]<=-137; ws[1][1 ][21]<=   9; ws[1][1 ][22]<= 103; ws[1][1 ][23]<=   4; ws[1][1 ][24]<=-171; ws[1][1 ][25]<=-191; ws[1][1 ][26]<=-114; ws[1][1 ][27]<=-134; ws[1][1 ][28]<= -27; ws[1][1 ][29]<=  55; ws[1][1 ][30]<= -56; ws[1][1 ][31]<=-208; ws[1][1 ][32]<=-237; ws[1][1 ][33]<=-142; ws[1][1 ][34]<= -70; ws[1][1 ][35]<=  34; ws[1][1 ][36]<=  37; ws[1][1 ][37]<=-133; ws[1][1 ][38]<=-246; ws[1][1 ][39]<=-119; ws[1][1 ][40]<= -66; ws[1][1 ][41]<= -46; ws[1][1 ][42]<=  97; ws[1][1 ][43]<=  53; ws[1][1 ][44]<=-123; ws[1][1 ][45]<=-159; ws[1][1 ][46]<=   8; ws[1][1 ][47]<=  81; ws[1][1 ][48]<=  19;
        ws[1][2 ][0]<= -67; ws[1][2 ][1]<=  17; ws[1][2 ][2]<= 105; ws[1][2 ][3]<= 139; ws[1][2 ][4]<= 109; ws[1][2 ][5]<=  62; ws[1][2 ][6]<= 123; ws[1][2 ][7]<= -86; ws[1][2 ][8]<= -64; ws[1][2 ][9]<=  22; ws[1][2 ][10]<=  73; ws[1][2 ][11]<=  92; ws[1][2 ][12]<=  75; ws[1][2 ][13]<= 165; ws[1][2 ][14]<=-109; ws[1][2 ][15]<=-102; ws[1][2 ][16]<= -13; ws[1][2 ][17]<=  48; ws[1][2 ][18]<=  56; ws[1][2 ][19]<=  48; ws[1][2 ][20]<= 148; ws[1][2 ][21]<=-115; ws[1][2 ][22]<=-177; ws[1][2 ][23]<= -52; ws[1][2 ][24]<= -22; ws[1][2 ][25]<=  52; ws[1][2 ][26]<=  77; ws[1][2 ][27]<= 167; ws[1][2 ][28]<=-125; ws[1][2 ][29]<=-202; ws[1][2 ][30]<= -59; ws[1][2 ][31]<=  21; ws[1][2 ][32]<=  59; ws[1][2 ][33]<=  91; ws[1][2 ][34]<= 156; ws[1][2 ][35]<=-188; ws[1][2 ][36]<=-115; ws[1][2 ][37]<=-107; ws[1][2 ][38]<= -13; ws[1][2 ][39]<=  67; ws[1][2 ][40]<=  93; ws[1][2 ][41]<= 153; ws[1][2 ][42]<=-160; ws[1][2 ][43]<=-166; ws[1][2 ][44]<= -55; ws[1][2 ][45]<= -39; ws[1][2 ][46]<=  35; ws[1][2 ][47]<= 110; ws[1][2 ][48]<= 215;
        ws[1][3 ][0]<=  12; ws[1][3 ][1]<=  64; ws[1][3 ][2]<=  92; ws[1][3 ][3]<=  94; ws[1][3 ][4]<=  -8; ws[1][3 ][5]<=-174; ws[1][3 ][6]<=-196; ws[1][3 ][7]<=  37; ws[1][3 ][8]<= 100; ws[1][3 ][9]<=  93; ws[1][3 ][10]<= 103; ws[1][3 ][11]<= -53; ws[1][3 ][12]<=-108; ws[1][3 ][13]<=-203; ws[1][3 ][14]<=  72; ws[1][3 ][15]<= 136; ws[1][3 ][16]<= 137; ws[1][3 ][17]<=  62; ws[1][3 ][18]<=  19; ws[1][3 ][19]<= -41; ws[1][3 ][20]<= -86; ws[1][3 ][21]<=  70; ws[1][3 ][22]<=  69; ws[1][3 ][23]<= 128; ws[1][3 ][24]<= 104; ws[1][3 ][25]<=  63; ws[1][3 ][26]<= -45; ws[1][3 ][27]<= -37; ws[1][3 ][28]<= -31; ws[1][3 ][29]<=  94; ws[1][3 ][30]<=  88; ws[1][3 ][31]<=  57; ws[1][3 ][32]<=  73; ws[1][3 ][33]<=   3; ws[1][3 ][34]<= -94; ws[1][3 ][35]<= -20; ws[1][3 ][36]<=  75; ws[1][3 ][37]<=  38; ws[1][3 ][38]<=  42; ws[1][3 ][39]<=  -3; ws[1][3 ][40]<= -64; ws[1][3 ][41]<= -91; ws[1][3 ][42]<= -87; ws[1][3 ][43]<=  -6; ws[1][3 ][44]<=  20; ws[1][3 ][45]<= -19; ws[1][3 ][46]<= -86; ws[1][3 ][47]<=-124; ws[1][3 ][48]<=-139;
        ws[1][4 ][0]<=  48; ws[1][4 ][1]<=  89; ws[1][4 ][2]<=  42; ws[1][4 ][3]<= -66; ws[1][4 ][4]<= -66; ws[1][4 ][5]<= -76; ws[1][4 ][6]<= -98; ws[1][4 ][7]<=  95; ws[1][4 ][8]<= 168; ws[1][4 ][9]<=  75; ws[1][4 ][10]<= -29; ws[1][4 ][11]<= -75; ws[1][4 ][12]<=   4; ws[1][4 ][13]<=-100; ws[1][4 ][14]<= 151; ws[1][4 ][15]<= 208; ws[1][4 ][16]<= 149; ws[1][4 ][17]<=  38; ws[1][4 ][18]<= -32; ws[1][4 ][19]<=  29; ws[1][4 ][20]<= -45; ws[1][4 ][21]<= 124; ws[1][4 ][22]<= 186; ws[1][4 ][23]<= 168; ws[1][4 ][24]<=   5; ws[1][4 ][25]<=  14; ws[1][4 ][26]<=  21; ws[1][4 ][27]<=  22; ws[1][4 ][28]<= 148; ws[1][4 ][29]<= 209; ws[1][4 ][30]<= 131; ws[1][4 ][31]<=   2; ws[1][4 ][32]<=  20; ws[1][4 ][33]<=   1; ws[1][4 ][34]<=  10; ws[1][4 ][35]<=  73; ws[1][4 ][36]<= 123; ws[1][4 ][37]<=  87; ws[1][4 ][38]<=   0; ws[1][4 ][39]<= -27; ws[1][4 ][40]<= -48; ws[1][4 ][41]<=  43; ws[1][4 ][42]<= 118; ws[1][4 ][43]<=  73; ws[1][4 ][44]<= 101; ws[1][4 ][45]<=   7; ws[1][4 ][46]<= -64; ws[1][4 ][47]<= -37; ws[1][4 ][48]<=   1;
        ws[1][5 ][0]<=-139; ws[1][5 ][1]<=-176; ws[1][5 ][2]<=-131; ws[1][5 ][3]<= -89; ws[1][5 ][4]<=-112; ws[1][5 ][5]<= -54; ws[1][5 ][6]<=  -3; ws[1][5 ][7]<=-117; ws[1][5 ][8]<=-168; ws[1][5 ][9]<=-112; ws[1][5 ][10]<= -95; ws[1][5 ][11]<= -87; ws[1][5 ][12]<=  17; ws[1][5 ][13]<=  78; ws[1][5 ][14]<=-101; ws[1][5 ][15]<=-163; ws[1][5 ][16]<=-122; ws[1][5 ][17]<= -74; ws[1][5 ][18]<=  15; ws[1][5 ][19]<=  34; ws[1][5 ][20]<=  76; ws[1][5 ][21]<= -29; ws[1][5 ][22]<=-151; ws[1][5 ][23]<= -80; ws[1][5 ][24]<=   1; ws[1][5 ][25]<=   4; ws[1][5 ][26]<=   3; ws[1][5 ][27]<=  50; ws[1][5 ][28]<=  14; ws[1][5 ][29]<=-100; ws[1][5 ][30]<= -29; ws[1][5 ][31]<=  18; ws[1][5 ][32]<=  37; ws[1][5 ][33]<=  51; ws[1][5 ][34]<= 149; ws[1][5 ][35]<=  17; ws[1][5 ][36]<= -44; ws[1][5 ][37]<=  35; ws[1][5 ][38]<=  55; ws[1][5 ][39]<= 129; ws[1][5 ][40]<= 133; ws[1][5 ][41]<= 206; ws[1][5 ][42]<=  61; ws[1][5 ][43]<= -35; ws[1][5 ][44]<=  25; ws[1][5 ][45]<= 102; ws[1][5 ][46]<= 109; ws[1][5 ][47]<= 207; ws[1][5 ][48]<= 257;
        ws[1][6 ][0]<= 146; ws[1][6 ][1]<= 168; ws[1][6 ][2]<=  60; ws[1][6 ][3]<= -26; ws[1][6 ][4]<=  29; ws[1][6 ][5]<=  11; ws[1][6 ][6]<=  14; ws[1][6 ][7]<= 167; ws[1][6 ][8]<=  90; ws[1][6 ][9]<=  56; ws[1][6 ][10]<=  25; ws[1][6 ][11]<=  33; ws[1][6 ][12]<=  20; ws[1][6 ][13]<=  93; ws[1][6 ][14]<=  97; ws[1][6 ][15]<= 129; ws[1][6 ][16]<=  13; ws[1][6 ][17]<=  18; ws[1][6 ][18]<= -35; ws[1][6 ][19]<=  -9; ws[1][6 ][20]<=  93; ws[1][6 ][21]<= 141; ws[1][6 ][22]<=  91; ws[1][6 ][23]<=  54; ws[1][6 ][24]<= -38; ws[1][6 ][25]<=  -2; ws[1][6 ][26]<=  36; ws[1][6 ][27]<=  56; ws[1][6 ][28]<= 153; ws[1][6 ][29]<= 129; ws[1][6 ][30]<=  75; ws[1][6 ][31]<=  -3; ws[1][6 ][32]<=   9; ws[1][6 ][33]<=  -3; ws[1][6 ][34]<=  40; ws[1][6 ][35]<= 143; ws[1][6 ][36]<= 157; ws[1][6 ][37]<= 105; ws[1][6 ][38]<=  77; ws[1][6 ][39]<=  35; ws[1][6 ][40]<=  69; ws[1][6 ][41]<=  81; ws[1][6 ][42]<= 204; ws[1][6 ][43]<= 187; ws[1][6 ][44]<=  89; ws[1][6 ][45]<=  82; ws[1][6 ][46]<=  56; ws[1][6 ][47]<=  81; ws[1][6 ][48]<=  60;
        ws[1][7 ][0]<=  20; ws[1][7 ][1]<=  54; ws[1][7 ][2]<= 160; ws[1][7 ][3]<= 182; ws[1][7 ][4]<= 133; ws[1][7 ][5]<=  82; ws[1][7 ][6]<= -26; ws[1][7 ][7]<= -19; ws[1][7 ][8]<=  52; ws[1][7 ][9]<= 231; ws[1][7 ][10]<= 202; ws[1][7 ][11]<=  67; ws[1][7 ][12]<=  40; ws[1][7 ][13]<= -47; ws[1][7 ][14]<= -37; ws[1][7 ][15]<= 104; ws[1][7 ][16]<= 219; ws[1][7 ][17]<= 137; ws[1][7 ][18]<=  80; ws[1][7 ][19]<= -34; ws[1][7 ][20]<= -30; ws[1][7 ][21]<=  56; ws[1][7 ][22]<= 175; ws[1][7 ][23]<= 183; ws[1][7 ][24]<=  81; ws[1][7 ][25]<=  -1; ws[1][7 ][26]<= -95; ws[1][7 ][27]<= -80; ws[1][7 ][28]<=  82; ws[1][7 ][29]<= 170; ws[1][7 ][30]<= 101; ws[1][7 ][31]<= -15; ws[1][7 ][32]<= -47; ws[1][7 ][33]<= -65; ws[1][7 ][34]<= -33; ws[1][7 ][35]<= 112; ws[1][7 ][36]<= 106; ws[1][7 ][37]<=  68; ws[1][7 ][38]<=  -3; ws[1][7 ][39]<=-113; ws[1][7 ][40]<=-121; ws[1][7 ][41]<= -57; ws[1][7 ][42]<=  31; ws[1][7 ][43]<=  95; ws[1][7 ][44]<=  40; ws[1][7 ][45]<= -20; ws[1][7 ][46]<=-130; ws[1][7 ][47]<= -85; ws[1][7 ][48]<= -89;
        ws[1][8 ][0]<=  64; ws[1][8 ][1]<= -59; ws[1][8 ][2]<= -60; ws[1][8 ][3]<=   9; ws[1][8 ][4]<=  43; ws[1][8 ][5]<=  43; ws[1][8 ][6]<= -20; ws[1][8 ][7]<=  66; ws[1][8 ][8]<= -38; ws[1][8 ][9]<= -52; ws[1][8 ][10]<= -54; ws[1][8 ][11]<=  36; ws[1][8 ][12]<=  90; ws[1][8 ][13]<=  18; ws[1][8 ][14]<=  28; ws[1][8 ][15]<= -23; ws[1][8 ][16]<=-105; ws[1][8 ][17]<= -15; ws[1][8 ][18]<= 137; ws[1][8 ][19]<= 155; ws[1][8 ][20]<=  61; ws[1][8 ][21]<=  27; ws[1][8 ][22]<= -60; ws[1][8 ][23]<= -64; ws[1][8 ][24]<= -35; ws[1][8 ][25]<= 148; ws[1][8 ][26]<= 121; ws[1][8 ][27]<=  76; ws[1][8 ][28]<=  35; ws[1][8 ][29]<=  35; ws[1][8 ][30]<=  -1; ws[1][8 ][31]<=  44; ws[1][8 ][32]<= 132; ws[1][8 ][33]<= 135; ws[1][8 ][34]<=  41; ws[1][8 ][35]<= 126; ws[1][8 ][36]<=  72; ws[1][8 ][37]<=  55; ws[1][8 ][38]<=  17; ws[1][8 ][39]<=  32; ws[1][8 ][40]<=  67; ws[1][8 ][41]<=  58; ws[1][8 ][42]<= 133; ws[1][8 ][43]<= 124; ws[1][8 ][44]<= 158; ws[1][8 ][45]<=  41; ws[1][8 ][46]<=  22; ws[1][8 ][47]<=  13; ws[1][8 ][48]<=  32;
        ws[1][9 ][0]<= -55; ws[1][9 ][1]<=  35; ws[1][9 ][2]<=  87; ws[1][9 ][3]<=  21; ws[1][9 ][4]<= -57; ws[1][9 ][5]<= -28; ws[1][9 ][6]<=  68; ws[1][9 ][7]<= -87; ws[1][9 ][8]<=-194; ws[1][9 ][9]<=-127; ws[1][9 ][10]<= -72; ws[1][9 ][11]<= -44; ws[1][9 ][12]<=   6; ws[1][9 ][13]<=  80; ws[1][9 ][14]<=-168; ws[1][9 ][15]<=-261; ws[1][9 ][16]<=-168; ws[1][9 ][17]<=  28; ws[1][9 ][18]<=  50; ws[1][9 ][19]<=  22; ws[1][9 ][20]<=  64; ws[1][9 ][21]<=-151; ws[1][9 ][22]<=-276; ws[1][9 ][23]<=-125; ws[1][9 ][24]<= 125; ws[1][9 ][25]<= 147; ws[1][9 ][26]<=  11; ws[1][9 ][27]<=  79; ws[1][9 ][28]<= -43; ws[1][9 ][29]<=-140; ws[1][9 ][30]<=  -3; ws[1][9 ][31]<= 181; ws[1][9 ][32]<= 138; ws[1][9 ][33]<=  -6; ws[1][9 ][34]<=   4; ws[1][9 ][35]<= -34; ws[1][9 ][36]<=  -8; ws[1][9 ][37]<=  73; ws[1][9 ][38]<= 218; ws[1][9 ][39]<= 159; ws[1][9 ][40]<=  46; ws[1][9 ][41]<=   1; ws[1][9 ][42]<=  -8; ws[1][9 ][43]<= -15; ws[1][9 ][44]<=  82; ws[1][9 ][45]<= 129; ws[1][9 ][46]<= 160; ws[1][9 ][47]<=  37; ws[1][9 ][48]<=  10;
        ws[1][10][0]<=  41; ws[1][10][1]<= -45; ws[1][10][2]<= -64; ws[1][10][3]<=   9; ws[1][10][4]<=  13; ws[1][10][5]<= -11; ws[1][10][6]<=  40; ws[1][10][7]<=  60; ws[1][10][8]<=  -8; ws[1][10][9]<=   2; ws[1][10][10]<=  17; ws[1][10][11]<=  79; ws[1][10][12]<=  26; ws[1][10][13]<=  37; ws[1][10][14]<=  21; ws[1][10][15]<=  12; ws[1][10][16]<=  39; ws[1][10][17]<=  63; ws[1][10][18]<=  99; ws[1][10][19]<=  83; ws[1][10][20]<=  45; ws[1][10][21]<=  41; ws[1][10][22]<=  50; ws[1][10][23]<=  77; ws[1][10][24]<= 152; ws[1][10][25]<= 142; ws[1][10][26]<=  39; ws[1][10][27]<=  53; ws[1][10][28]<=  81; ws[1][10][29]<=  45; ws[1][10][30]<=  47; ws[1][10][31]<= 174; ws[1][10][32]<= 160; ws[1][10][33]<=  71; ws[1][10][34]<=  65; ws[1][10][35]<=  78; ws[1][10][36]<=  47; ws[1][10][37]<= 104; ws[1][10][38]<= 165; ws[1][10][39]<= 107; ws[1][10][40]<= 111; ws[1][10][41]<=  86; ws[1][10][42]<=  48; ws[1][10][43]<=  55; ws[1][10][44]<=  62; ws[1][10][45]<= 113; ws[1][10][46]<= 170; ws[1][10][47]<= 142; ws[1][10][48]<=  53;
        ws[1][11][0]<=  74; ws[1][11][1]<= -55; ws[1][11][2]<= -47; ws[1][11][3]<= -22; ws[1][11][4]<=  -2; ws[1][11][5]<=  -1; ws[1][11][6]<= -59; ws[1][11][7]<= -67; ws[1][11][8]<= -52; ws[1][11][9]<= -29; ws[1][11][10]<=  -9; ws[1][11][11]<=  -8; ws[1][11][12]<=  -9; ws[1][11][13]<=  10; ws[1][11][14]<=-116; ws[1][11][15]<=-138; ws[1][11][16]<=-119; ws[1][11][17]<= -50; ws[1][11][18]<= -37; ws[1][11][19]<= -18; ws[1][11][20]<= -10; ws[1][11][21]<=-122; ws[1][11][22]<=-186; ws[1][11][23]<=-155; ws[1][11][24]<= -67; ws[1][11][25]<= -57; ws[1][11][26]<=  -2; ws[1][11][27]<=  17; ws[1][11][28]<= -76; ws[1][11][29]<=-108; ws[1][11][30]<=-139; ws[1][11][31]<= -82; ws[1][11][32]<=  -3; ws[1][11][33]<=  10; ws[1][11][34]<=  73; ws[1][11][35]<= -11; ws[1][11][36]<= -78; ws[1][11][37]<=-141; ws[1][11][38]<=-100; ws[1][11][39]<= -14; ws[1][11][40]<=  42; ws[1][11][41]<=  91; ws[1][11][42]<= -68; ws[1][11][43]<= -86; ws[1][11][44]<= -82; ws[1][11][45]<= -60; ws[1][11][46]<=  28; ws[1][11][47]<= 154; ws[1][11][48]<= 154;
        ws[1][12][0]<=   7; ws[1][12][1]<=-140; ws[1][12][2]<=-230; ws[1][12][3]<=-136; ws[1][12][4]<= -99; ws[1][12][5]<=   2; ws[1][12][6]<= -93; ws[1][12][7]<=   6; ws[1][12][8]<=-116; ws[1][12][9]<=-198; ws[1][12][10]<=-105; ws[1][12][11]<= -75; ws[1][12][12]<= -15; ws[1][12][13]<= -16; ws[1][12][14]<= -26; ws[1][12][15]<=-118; ws[1][12][16]<=-138; ws[1][12][17]<=-101; ws[1][12][18]<=  -4; ws[1][12][19]<=  -6; ws[1][12][20]<=  25; ws[1][12][21]<=   7; ws[1][12][22]<= -51; ws[1][12][23]<=-113; ws[1][12][24]<=-118; ws[1][12][25]<= -55; ws[1][12][26]<=  16; ws[1][12][27]<=  36; ws[1][12][28]<=  34; ws[1][12][29]<= -37; ws[1][12][30]<=-130; ws[1][12][31]<=-127; ws[1][12][32]<= -56; ws[1][12][33]<=  58; ws[1][12][34]<=  36; ws[1][12][35]<=  61; ws[1][12][36]<=   5; ws[1][12][37]<= -90; ws[1][12][38]<= -38; ws[1][12][39]<=  18; ws[1][12][40]<=  56; ws[1][12][41]<=  51; ws[1][12][42]<=  83; ws[1][12][43]<=  27; ws[1][12][44]<=   1; ws[1][12][45]<= -26; ws[1][12][46]<= -29; ws[1][12][47]<=  38; ws[1][12][48]<=  47;
        ws[1][13][0]<=-135; ws[1][13][1]<= -96; ws[1][13][2]<=-143; ws[1][13][3]<=-115; ws[1][13][4]<= -98; ws[1][13][5]<= -35; ws[1][13][6]<=  30; ws[1][13][7]<=-156; ws[1][13][8]<=-174; ws[1][13][9]<=-132; ws[1][13][10]<=-117; ws[1][13][11]<= -74; ws[1][13][12]<=  -9; ws[1][13][13]<=  49; ws[1][13][14]<=-130; ws[1][13][15]<=-157; ws[1][13][16]<=-186; ws[1][13][17]<= -66; ws[1][13][18]<=  40; ws[1][13][19]<=  39; ws[1][13][20]<=  59; ws[1][13][21]<= -93; ws[1][13][22]<=-152; ws[1][13][23]<= -55; ws[1][13][24]<=  53; ws[1][13][25]<= 129; ws[1][13][26]<=  67; ws[1][13][27]<=  75; ws[1][13][28]<=  -9; ws[1][13][29]<= -28; ws[1][13][30]<=  19; ws[1][13][31]<= 103; ws[1][13][32]<= 180; ws[1][13][33]<= 106; ws[1][13][34]<=  70; ws[1][13][35]<=  -1; ws[1][13][36]<= -27; ws[1][13][37]<= 107; ws[1][13][38]<= 176; ws[1][13][39]<= 173; ws[1][13][40]<=  67; ws[1][13][41]<=  87; ws[1][13][42]<=  -8; ws[1][13][43]<= -85; ws[1][13][44]<= 117; ws[1][13][45]<= 160; ws[1][13][46]<= 103; ws[1][13][47]<=  73; ws[1][13][48]<=  44;
        ws[1][14][0]<= -61; ws[1][14][1]<= -63; ws[1][14][2]<=-113; ws[1][14][3]<=-138; ws[1][14][4]<= -45; ws[1][14][5]<= -16; ws[1][14][6]<=  19; ws[1][14][7]<= -75; ws[1][14][8]<=  -4; ws[1][14][9]<= -96; ws[1][14][10]<=-150; ws[1][14][11]<=-118; ws[1][14][12]<= -46; ws[1][14][13]<= -23; ws[1][14][14]<=  22; ws[1][14][15]<=  78; ws[1][14][16]<= -90; ws[1][14][17]<=-173; ws[1][14][18]<=-156; ws[1][14][19]<= -17; ws[1][14][20]<=-102; ws[1][14][21]<=  93; ws[1][14][22]<= 117; ws[1][14][23]<=  37; ws[1][14][24]<=-146; ws[1][14][25]<= -88; ws[1][14][26]<= -71; ws[1][14][27]<= -85; ws[1][14][28]<= 114; ws[1][14][29]<= 171; ws[1][14][30]<=  -3; ws[1][14][31]<= -55; ws[1][14][32]<=-104; ws[1][14][33]<= -60; ws[1][14][34]<= -49; ws[1][14][35]<= 162; ws[1][14][36]<= 190; ws[1][14][37]<=  19; ws[1][14][38]<= -88; ws[1][14][39]<=-112; ws[1][14][40]<= -73; ws[1][14][41]<= -96; ws[1][14][42]<= 186; ws[1][14][43]<= 149; ws[1][14][44]<= 116; ws[1][14][45]<= -87; ws[1][14][46]<=-106; ws[1][14][47]<=   4; ws[1][14][48]<= -83;
        ws[1][15][0]<=  96; ws[1][15][1]<= -20; ws[1][15][2]<=-106; ws[1][15][3]<= -38; ws[1][15][4]<= 166; ws[1][15][5]<= 290; ws[1][15][6]<= 285; ws[1][15][7]<=   4; ws[1][15][8]<=  -1; ws[1][15][9]<= -28; ws[1][15][10]<=  -7; ws[1][15][11]<=  84; ws[1][15][12]<= 176; ws[1][15][13]<= 181; ws[1][15][14]<= -43; ws[1][15][15]<= -28; ws[1][15][16]<=  54; ws[1][15][17]<=  29; ws[1][15][18]<= -10; ws[1][15][19]<=  35; ws[1][15][20]<=  88; ws[1][15][21]<= -34; ws[1][15][22]<=  50; ws[1][15][23]<= 116; ws[1][15][24]<= -67; ws[1][15][25]<=-131; ws[1][15][26]<= -92; ws[1][15][27]<= -35; ws[1][15][28]<= -44; ws[1][15][29]<=  39; ws[1][15][30]<=  88; ws[1][15][31]<= -96; ws[1][15][32]<=-249; ws[1][15][33]<=-124; ws[1][15][34]<= -73; ws[1][15][35]<=  19; ws[1][15][36]<=  12; ws[1][15][37]<= 121; ws[1][15][38]<= -40; ws[1][15][39]<=-222; ws[1][15][40]<=-200; ws[1][15][41]<=-127; ws[1][15][42]<=  -2; ws[1][15][43]<= -40; ws[1][15][44]<=  22; ws[1][15][45]<=   2; ws[1][15][46]<=-175; ws[1][15][47]<=-170; ws[1][15][48]<=-164;

        ws[2][0 ][0]<=  79; ws[2][0 ][1]<= -24; ws[2][0 ][2]<= -43; ws[2][0 ][3]<= -57; ws[2][0 ][4]<= -64; ws[2][0 ][5]<=  22; ws[2][0 ][6]<= 130; ws[2][0 ][7]<=  -8; ws[2][0 ][8]<= -10; ws[2][0 ][9]<= -52; ws[2][0 ][10]<=-117; ws[2][0 ][11]<= -43; ws[2][0 ][12]<=  85; ws[2][0 ][13]<=  95; ws[2][0 ][14]<= -49; ws[2][0 ][15]<= -87; ws[2][0 ][16]<=-132; ws[2][0 ][17]<= -82; ws[2][0 ][18]<=  10; ws[2][0 ][19]<=  44; ws[2][0 ][20]<= 200; ws[2][0 ][21]<= -22; ws[2][0 ][22]<= -37; ws[2][0 ][23]<=-109; ws[2][0 ][24]<=-130; ws[2][0 ][25]<=  11; ws[2][0 ][26]<= 150; ws[2][0 ][27]<= 216; ws[2][0 ][28]<= -23; ws[2][0 ][29]<= -63; ws[2][0 ][30]<=-108; ws[2][0 ][31]<= -36; ws[2][0 ][32]<=   7; ws[2][0 ][33]<= 109; ws[2][0 ][34]<= 269; ws[2][0 ][35]<= -42; ws[2][0 ][36]<=  -2; ws[2][0 ][37]<= -39; ws[2][0 ][38]<= -12; ws[2][0 ][39]<=  -2; ws[2][0 ][40]<= 147; ws[2][0 ][41]<= 286; ws[2][0 ][42]<= -31; ws[2][0 ][43]<=  25; ws[2][0 ][44]<=  63; ws[2][0 ][45]<=  78; ws[2][0 ][46]<=  97; ws[2][0 ][47]<= 158; ws[2][0 ][48]<= 306;
        ws[2][1 ][0]<= -95; ws[2][1 ][1]<= -42; ws[2][1 ][2]<= -79; ws[2][1 ][3]<=-189; ws[2][1 ][4]<=-193; ws[2][1 ][5]<= -17; ws[2][1 ][6]<=  88; ws[2][1 ][7]<= -99; ws[2][1 ][8]<= -36; ws[2][1 ][9]<= -18; ws[2][1 ][10]<=-115; ws[2][1 ][11]<=-129; ws[2][1 ][12]<= -27; ws[2][1 ][13]<= -11; ws[2][1 ][14]<=-122; ws[2][1 ][15]<= -51; ws[2][1 ][16]<=  23; ws[2][1 ][17]<= -21; ws[2][1 ][18]<=-125; ws[2][1 ][19]<= -60; ws[2][1 ][20]<=  -3; ws[2][1 ][21]<= -15; ws[2][1 ][22]<=  -7; ws[2][1 ][23]<=  10; ws[2][1 ][24]<=  17; ws[2][1 ][25]<=-137; ws[2][1 ][26]<=-131; ws[2][1 ][27]<= -74; ws[2][1 ][28]<= -15; ws[2][1 ][29]<=  69; ws[2][1 ][30]<=   4; ws[2][1 ][31]<= -25; ws[2][1 ][32]<=-113; ws[2][1 ][33]<=-170; ws[2][1 ][34]<=-133; ws[2][1 ][35]<= -49; ws[2][1 ][36]<= -31; ws[2][1 ][37]<= -61; ws[2][1 ][38]<= -81; ws[2][1 ][39]<= -81; ws[2][1 ][40]<=-129; ws[2][1 ][41]<=-128; ws[2][1 ][42]<=-211; ws[2][1 ][43]<=-153; ws[2][1 ][44]<=-183; ws[2][1 ][45]<=-134; ws[2][1 ][46]<= -48; ws[2][1 ][47]<=-135; ws[2][1 ][48]<=-139;
        ws[2][2 ][0]<=  87; ws[2][2 ][1]<=-172; ws[2][2 ][2]<=-175; ws[2][2 ][3]<=  90; ws[2][2 ][4]<= 187; ws[2][2 ][5]<= 134; ws[2][2 ][6]<= 121; ws[2][2 ][7]<=  75; ws[2][2 ][8]<= -69; ws[2][2 ][9]<=-128; ws[2][2 ][10]<=  68; ws[2][2 ][11]<= 215; ws[2][2 ][12]<= 162; ws[2][2 ][13]<=  96; ws[2][2 ][14]<=  73; ws[2][2 ][15]<= -29; ws[2][2 ][16]<=-116; ws[2][2 ][17]<=  44; ws[2][2 ][18]<= 160; ws[2][2 ][19]<= 109; ws[2][2 ][20]<= 117; ws[2][2 ][21]<=  72; ws[2][2 ][22]<= -52; ws[2][2 ][23]<=-118; ws[2][2 ][24]<= -44; ws[2][2 ][25]<=  91; ws[2][2 ][26]<=  66; ws[2][2 ][27]<=  80; ws[2][2 ][28]<=  26; ws[2][2 ][29]<= -17; ws[2][2 ][30]<=-206; ws[2][2 ][31]<=-160; ws[2][2 ][32]<= -35; ws[2][2 ][33]<= -16; ws[2][2 ][34]<= -66; ws[2][2 ][35]<= -13; ws[2][2 ][36]<=  40; ws[2][2 ][37]<=-169; ws[2][2 ][38]<=-202; ws[2][2 ][39]<=-118; ws[2][2 ][40]<= -25; ws[2][2 ][41]<=-170; ws[2][2 ][42]<= -21; ws[2][2 ][43]<=  63; ws[2][2 ][44]<= -48; ws[2][2 ][45]<= -97; ws[2][2 ][46]<= -20; ws[2][2 ][47]<= -57; ws[2][2 ][48]<=-223;
        ws[2][3 ][0]<=  96; ws[2][3 ][1]<=  60; ws[2][3 ][2]<= -27; ws[2][3 ][3]<=  23; ws[2][3 ][4]<= -57; ws[2][3 ][5]<=-221; ws[2][3 ][6]<=-162; ws[2][3 ][7]<= -18; ws[2][3 ][8]<= -24; ws[2][3 ][9]<= -27; ws[2][3 ][10]<=  72; ws[2][3 ][11]<= 106; ws[2][3 ][12]<= -14; ws[2][3 ][13]<=  -5; ws[2][3 ][14]<=  12; ws[2][3 ][15]<= -55; ws[2][3 ][16]<=   2; ws[2][3 ][17]<= 211; ws[2][3 ][18]<= 257; ws[2][3 ][19]<= 173; ws[2][3 ][20]<=  22; ws[2][3 ][21]<= -15; ws[2][3 ][22]<=  25; ws[2][3 ][23]<=   5; ws[2][3 ][24]<= 251; ws[2][3 ][25]<= 331; ws[2][3 ][26]<= 172; ws[2][3 ][27]<= -32; ws[2][3 ][28]<=  41; ws[2][3 ][29]<=  -1; ws[2][3 ][30]<=  23; ws[2][3 ][31]<=  91; ws[2][3 ][32]<= 266; ws[2][3 ][33]<= 104; ws[2][3 ][34]<=-121; ws[2][3 ][35]<= -80; ws[2][3 ][36]<=  38; ws[2][3 ][37]<= -24; ws[2][3 ][38]<= -19; ws[2][3 ][39]<= 110; ws[2][3 ][40]<=  99; ws[2][3 ][41]<=-104; ws[2][3 ][42]<=-147; ws[2][3 ][43]<=  24; ws[2][3 ][44]<=   3; ws[2][3 ][45]<= -85; ws[2][3 ][46]<= -49; ws[2][3 ][47]<=  89; ws[2][3 ][48]<= -44;
        ws[2][4 ][0]<=  87; ws[2][4 ][1]<= 185; ws[2][4 ][2]<= 130; ws[2][4 ][3]<=  32; ws[2][4 ][4]<=   3; ws[2][4 ][5]<=  71; ws[2][4 ][6]<=  12; ws[2][4 ][7]<= 155; ws[2][4 ][8]<= 140; ws[2][4 ][9]<= 112; ws[2][4 ][10]<=  76; ws[2][4 ][11]<=  27; ws[2][4 ][12]<=  55; ws[2][4 ][13]<=  21; ws[2][4 ][14]<= 114; ws[2][4 ][15]<= 196; ws[2][4 ][16]<=  61; ws[2][4 ][17]<=  -1; ws[2][4 ][18]<=  39; ws[2][4 ][19]<=  43; ws[2][4 ][20]<=  59; ws[2][4 ][21]<=  82; ws[2][4 ][22]<= 144; ws[2][4 ][23]<= 103; ws[2][4 ][24]<=  -4; ws[2][4 ][25]<= -15; ws[2][4 ][26]<=   9; ws[2][4 ][27]<=  33; ws[2][4 ][28]<=  85; ws[2][4 ][29]<= 182; ws[2][4 ][30]<=  94; ws[2][4 ][31]<=  11; ws[2][4 ][32]<=  30; ws[2][4 ][33]<=  66; ws[2][4 ][34]<=   6; ws[2][4 ][35]<= 130; ws[2][4 ][36]<= 195; ws[2][4 ][37]<= 112; ws[2][4 ][38]<=   1; ws[2][4 ][39]<=  15; ws[2][4 ][40]<=  50; ws[2][4 ][41]<=  35; ws[2][4 ][42]<= 123; ws[2][4 ][43]<= 163; ws[2][4 ][44]<= 122; ws[2][4 ][45]<=  31; ws[2][4 ][46]<=  33; ws[2][4 ][47]<=  79; ws[2][4 ][48]<=  80;
        ws[2][5 ][0]<=-106; ws[2][5 ][1]<=  25; ws[2][5 ][2]<=  66; ws[2][5 ][3]<= 109; ws[2][5 ][4]<=  43; ws[2][5 ][5]<=-108; ws[2][5 ][6]<=-117; ws[2][5 ][7]<= -78; ws[2][5 ][8]<=  62; ws[2][5 ][9]<=  87; ws[2][5 ][10]<= 106; ws[2][5 ][11]<=   1; ws[2][5 ][12]<= -22; ws[2][5 ][13]<=-161; ws[2][5 ][14]<= -14; ws[2][5 ][15]<=  26; ws[2][5 ][16]<= -24; ws[2][5 ][17]<=  17; ws[2][5 ][18]<=  87; ws[2][5 ][19]<= -55; ws[2][5 ][20]<=-143; ws[2][5 ][21]<= -82; ws[2][5 ][22]<=  -9; ws[2][5 ][23]<= -68; ws[2][5 ][24]<= -35; ws[2][5 ][25]<=  26; ws[2][5 ][26]<= -34; ws[2][5 ][27]<=-115; ws[2][5 ][28]<= -47; ws[2][5 ][29]<= -70; ws[2][5 ][30]<=-126; ws[2][5 ][31]<=-141; ws[2][5 ][32]<= -23; ws[2][5 ][33]<= -30; ws[2][5 ][34]<= -87; ws[2][5 ][35]<= -24; ws[2][5 ][36]<= -42; ws[2][5 ][37]<=-148; ws[2][5 ][38]<=-209; ws[2][5 ][39]<= -56; ws[2][5 ][40]<= -18; ws[2][5 ][41]<= -49; ws[2][5 ][42]<= 111; ws[2][5 ][43]<=  44; ws[2][5 ][44]<=-163; ws[2][5 ][45]<=-237; ws[2][5 ][46]<= -50; ws[2][5 ][47]<=  17; ws[2][5 ][48]<= -90;
        ws[2][6 ][0]<= -68; ws[2][6 ][1]<=-106; ws[2][6 ][2]<=-123; ws[2][6 ][3]<= -78; ws[2][6 ][4]<=  86; ws[2][6 ][5]<= 136; ws[2][6 ][6]<= 126; ws[2][6 ][7]<= -29; ws[2][6 ][8]<= -72; ws[2][6 ][9]<=-155; ws[2][6 ][10]<= -87; ws[2][6 ][11]<=  72; ws[2][6 ][12]<= 164; ws[2][6 ][13]<= 174; ws[2][6 ][14]<=  87; ws[2][6 ][15]<= -32; ws[2][6 ][16]<=-154; ws[2][6 ][17]<=-121; ws[2][6 ][18]<=  27; ws[2][6 ][19]<= 166; ws[2][6 ][20]<= 161; ws[2][6 ][21]<=  57; ws[2][6 ][22]<= -76; ws[2][6 ][23]<=-172; ws[2][6 ][24]<=-163; ws[2][6 ][25]<=  26; ws[2][6 ][26]<= 125; ws[2][6 ][27]<= 168; ws[2][6 ][28]<= -28; ws[2][6 ][29]<= -30; ws[2][6 ][30]<=-135; ws[2][6 ][31]<= -85; ws[2][6 ][32]<= -16; ws[2][6 ][33]<= 107; ws[2][6 ][34]<= 143; ws[2][6 ][35]<=-104; ws[2][6 ][36]<= -32; ws[2][6 ][37]<= -29; ws[2][6 ][38]<= -12; ws[2][6 ][39]<= -34; ws[2][6 ][40]<=  53; ws[2][6 ][41]<= 164; ws[2][6 ][42]<=-153; ws[2][6 ][43]<= -54; ws[2][6 ][44]<=   2; ws[2][6 ][45]<=  40; ws[2][6 ][46]<=  66; ws[2][6 ][47]<= 137; ws[2][6 ][48]<= 195;
        ws[2][7 ][0]<=  53; ws[2][7 ][1]<=  25; ws[2][7 ][2]<=  40; ws[2][7 ][3]<=   5; ws[2][7 ][4]<=  -3; ws[2][7 ][5]<=-164; ws[2][7 ][6]<=-162; ws[2][7 ][7]<=  60; ws[2][7 ][8]<=  29; ws[2][7 ][9]<= -23; ws[2][7 ][10]<=   4; ws[2][7 ][11]<= -25; ws[2][7 ][12]<=  -1; ws[2][7 ][13]<= -83; ws[2][7 ][14]<=  46; ws[2][7 ][15]<= -17; ws[2][7 ][16]<=   7; ws[2][7 ][17]<=  55; ws[2][7 ][18]<= 104; ws[2][7 ][19]<=  87; ws[2][7 ][20]<=  56; ws[2][7 ][21]<=  97; ws[2][7 ][22]<=  21; ws[2][7 ][23]<=  50; ws[2][7 ][24]<= 164; ws[2][7 ][25]<= 217; ws[2][7 ][26]<= 142; ws[2][7 ][27]<=   9; ws[2][7 ][28]<=  72; ws[2][7 ][29]<=  82; ws[2][7 ][30]<= 160; ws[2][7 ][31]<= 249; ws[2][7 ][32]<= 249; ws[2][7 ][33]<= 115; ws[2][7 ][34]<=  69; ws[2][7 ][35]<=  70; ws[2][7 ][36]<=  37; ws[2][7 ][37]<=  91; ws[2][7 ][38]<= 170; ws[2][7 ][39]<= 173; ws[2][7 ][40]<=  76; ws[2][7 ][41]<=  77; ws[2][7 ][42]<= -77; ws[2][7 ][43]<=-136; ws[2][7 ][44]<= -24; ws[2][7 ][45]<=  75; ws[2][7 ][46]<=  82; ws[2][7 ][47]<= 111; ws[2][7 ][48]<=  33;
        ws[2][8 ][0]<=   6; ws[2][8 ][1]<= -25; ws[2][8 ][2]<=  83; ws[2][8 ][3]<= 132; ws[2][8 ][4]<= 108; ws[2][8 ][5]<=  37; ws[2][8 ][6]<= 109; ws[2][8 ][7]<=  11; ws[2][8 ][8]<= -14; ws[2][8 ][9]<=  81; ws[2][8 ][10]<= 139; ws[2][8 ][11]<= 132; ws[2][8 ][12]<=  81; ws[2][8 ][13]<=  68; ws[2][8 ][14]<=  93; ws[2][8 ][15]<=  39; ws[2][8 ][16]<=  40; ws[2][8 ][17]<=  96; ws[2][8 ][18]<= 146; ws[2][8 ][19]<= 132; ws[2][8 ][20]<=  68; ws[2][8 ][21]<= 112; ws[2][8 ][22]<=  -3; ws[2][8 ][23]<=  -4; ws[2][8 ][24]<= 114; ws[2][8 ][25]<= 184; ws[2][8 ][26]<= 154; ws[2][8 ][27]<=  97; ws[2][8 ][28]<=  28; ws[2][8 ][29]<= -32; ws[2][8 ][30]<=-100; ws[2][8 ][31]<=  15; ws[2][8 ][32]<=  95; ws[2][8 ][33]<= 164; ws[2][8 ][34]<=  47; ws[2][8 ][35]<= -39; ws[2][8 ][36]<= -75; ws[2][8 ][37]<=-153; ws[2][8 ][38]<= -32; ws[2][8 ][39]<=  72; ws[2][8 ][40]<=  81; ws[2][8 ][41]<=  10; ws[2][8 ][42]<=-112; ws[2][8 ][43]<= -88; ws[2][8 ][44]<= -59; ws[2][8 ][45]<=  -7; ws[2][8 ][46]<=  33; ws[2][8 ][47]<=   7; ws[2][8 ][48]<=   3;
        ws[2][9 ][0]<= -20; ws[2][9 ][1]<= -73; ws[2][9 ][2]<= -47; ws[2][9 ][3]<= -65; ws[2][9 ][4]<= -24; ws[2][9 ][5]<=  11; ws[2][9 ][6]<= -15; ws[2][9 ][7]<= -53; ws[2][9 ][8]<= -12; ws[2][9 ][9]<= -53; ws[2][9 ][10]<=  -9; ws[2][9 ][11]<= -27; ws[2][9 ][12]<= -28; ws[2][9 ][13]<=   5; ws[2][9 ][14]<= -80; ws[2][9 ][15]<= -87; ws[2][9 ][16]<= -50; ws[2][9 ][17]<= -62; ws[2][9 ][18]<= -42; ws[2][9 ][19]<= -66; ws[2][9 ][20]<= -49; ws[2][9 ][21]<= -41; ws[2][9 ][22]<= -80; ws[2][9 ][23]<= -68; ws[2][9 ][24]<= -28; ws[2][9 ][25]<= -46; ws[2][9 ][26]<= -72; ws[2][9 ][27]<= -71; ws[2][9 ][28]<= -82; ws[2][9 ][29]<= -36; ws[2][9 ][30]<= -56; ws[2][9 ][31]<= -85; ws[2][9 ][32]<=  -3; ws[2][9 ][33]<= -54; ws[2][9 ][34]<= -55; ws[2][9 ][35]<=-118; ws[2][9 ][36]<= -57; ws[2][9 ][37]<= -65; ws[2][9 ][38]<= -92; ws[2][9 ][39]<= -71; ws[2][9 ][40]<= -68; ws[2][9 ][41]<= -28; ws[2][9 ][42]<= -63; ws[2][9 ][43]<= -53; ws[2][9 ][44]<= -50; ws[2][9 ][45]<= -95; ws[2][9 ][46]<= -40; ws[2][9 ][47]<= -27; ws[2][9 ][48]<= -25;
        ws[2][10][0]<=-161; ws[2][10][1]<= -83; ws[2][10][2]<= -33; ws[2][10][3]<= -20; ws[2][10][4]<=-114; ws[2][10][5]<= -27; ws[2][10][6]<= -34; ws[2][10][7]<= -99; ws[2][10][8]<= -21; ws[2][10][9]<= -11; ws[2][10][10]<=   9; ws[2][10][11]<=  -6; ws[2][10][12]<= -36; ws[2][10][13]<= -25; ws[2][10][14]<=   7; ws[2][10][15]<=  98; ws[2][10][16]<=  45; ws[2][10][17]<=  30; ws[2][10][18]<=  18; ws[2][10][19]<=  40; ws[2][10][20]<=  51; ws[2][10][21]<=  76; ws[2][10][22]<=  88; ws[2][10][23]<=  99; ws[2][10][24]<= -19; ws[2][10][25]<= -30; ws[2][10][26]<=  50; ws[2][10][27]<=  36; ws[2][10][28]<=  63; ws[2][10][29]<=  77; ws[2][10][30]<=  28; ws[2][10][31]<=  41; ws[2][10][32]<=  -6; ws[2][10][33]<=  45; ws[2][10][34]<=  67; ws[2][10][35]<=  57; ws[2][10][36]<=  32; ws[2][10][37]<=  88; ws[2][10][38]<=  93; ws[2][10][39]<=  67; ws[2][10][40]<= 119; ws[2][10][41]<= 105; ws[2][10][42]<=  21; ws[2][10][43]<=  32; ws[2][10][44]<= 108; ws[2][10][45]<= 191; ws[2][10][46]<= 159; ws[2][10][47]<= 201; ws[2][10][48]<= 175;
        ws[2][11][0]<= 136; ws[2][11][1]<=-100; ws[2][11][2]<= -79; ws[2][11][3]<= -24; ws[2][11][4]<= -55; ws[2][11][5]<=  -2; ws[2][11][6]<=  49; ws[2][11][7]<=  82; ws[2][11][8]<= -81; ws[2][11][9]<= -31; ws[2][11][10]<= -69; ws[2][11][11]<= -19; ws[2][11][12]<=  24; ws[2][11][13]<=  59; ws[2][11][14]<=   3; ws[2][11][15]<=   3; ws[2][11][16]<=  -3; ws[2][11][17]<= -27; ws[2][11][18]<= -37; ws[2][11][19]<=  40; ws[2][11][20]<=  84; ws[2][11][21]<= -86; ws[2][11][22]<= -70; ws[2][11][23]<= -80; ws[2][11][24]<= -28; ws[2][11][25]<=  -6; ws[2][11][26]<=  64; ws[2][11][27]<= 131; ws[2][11][28]<=-112; ws[2][11][29]<= -88; ws[2][11][30]<=-135; ws[2][11][31]<=-163; ws[2][11][32]<= -99; ws[2][11][33]<=  39; ws[2][11][34]<=  27; ws[2][11][35]<=-131; ws[2][11][36]<= -74; ws[2][11][37]<=-156; ws[2][11][38]<=-174; ws[2][11][39]<=-180; ws[2][11][40]<= -39; ws[2][11][41]<= -39; ws[2][11][42]<= -62; ws[2][11][43]<= -36; ws[2][11][44]<=-104; ws[2][11][45]<=-153; ws[2][11][46]<= -88; ws[2][11][47]<= -50; ws[2][11][48]<= -84;
        ws[2][12][0]<= 108; ws[2][12][1]<=   8; ws[2][12][2]<=  15; ws[2][12][3]<=  55; ws[2][12][4]<=  16; ws[2][12][5]<=  76; ws[2][12][6]<=  55; ws[2][12][7]<= 139; ws[2][12][8]<=  93; ws[2][12][9]<=  39; ws[2][12][10]<= -50; ws[2][12][11]<= -71; ws[2][12][12]<=  18; ws[2][12][13]<=  69; ws[2][12][14]<=  48; ws[2][12][15]<= -24; ws[2][12][16]<= -66; ws[2][12][17]<=-121; ws[2][12][18]<=-148; ws[2][12][19]<= -17; ws[2][12][20]<= 104; ws[2][12][21]<= -37; ws[2][12][22]<= -32; ws[2][12][23]<=-176; ws[2][12][24]<=-194; ws[2][12][25]<=-134; ws[2][12][26]<= -14; ws[2][12][27]<=   1; ws[2][12][28]<= -98; ws[2][12][29]<= -78; ws[2][12][30]<=-183; ws[2][12][31]<=-107; ws[2][12][32]<= -98; ws[2][12][33]<= -65; ws[2][12][34]<= -64; ws[2][12][35]<= -96; ws[2][12][36]<=-141; ws[2][12][37]<= -65; ws[2][12][38]<= -45; ws[2][12][39]<= -22; ws[2][12][40]<= -37; ws[2][12][41]<=-145; ws[2][12][42]<= -48; ws[2][12][43]<=-132; ws[2][12][44]<= -77; ws[2][12][45]<=  41; ws[2][12][46]<=  10; ws[2][12][47]<= -69; ws[2][12][48]<=-222;
        ws[2][13][0]<= -67; ws[2][13][1]<= -88; ws[2][13][2]<=  15; ws[2][13][3]<= 107; ws[2][13][4]<= 105; ws[2][13][5]<=  -6; ws[2][13][6]<= -55; ws[2][13][7]<=-133; ws[2][13][8]<= -86; ws[2][13][9]<=  16; ws[2][13][10]<= 141; ws[2][13][11]<= 102; ws[2][13][12]<=  27; ws[2][13][13]<= -16; ws[2][13][14]<= -43; ws[2][13][15]<=-123; ws[2][13][16]<= -31; ws[2][13][17]<=  77; ws[2][13][18]<= 118; ws[2][13][19]<=  41; ws[2][13][20]<= -82; ws[2][13][21]<=  36; ws[2][13][22]<= -72; ws[2][13][23]<=  19; ws[2][13][24]<= 133; ws[2][13][25]<=  82; ws[2][13][26]<= -39; ws[2][13][27]<= -61; ws[2][13][28]<=  36; ws[2][13][29]<=  19; ws[2][13][30]<=  65; ws[2][13][31]<= 107; ws[2][13][32]<= 106; ws[2][13][33]<=  12; ws[2][13][34]<= -20; ws[2][13][35]<= 166; ws[2][13][36]<=  33; ws[2][13][37]<= 106; ws[2][13][38]<=  71; ws[2][13][39]<= 102; ws[2][13][40]<= 110; ws[2][13][41]<= -22; ws[2][13][42]<= 129; ws[2][13][43]<= 120; ws[2][13][44]<= 187; ws[2][13][45]<= 157; ws[2][13][46]<= 148; ws[2][13][47]<= 117; ws[2][13][48]<=  16;
        ws[2][14][0]<=  54; ws[2][14][1]<=  74; ws[2][14][2]<=  42; ws[2][14][3]<=   5; ws[2][14][4]<= -41; ws[2][14][5]<= -21; ws[2][14][6]<= -17; ws[2][14][7]<= -10; ws[2][14][8]<= -54; ws[2][14][9]<= -65; ws[2][14][10]<= -57; ws[2][14][11]<= -13; ws[2][14][12]<=  64; ws[2][14][13]<=  68; ws[2][14][14]<= -65; ws[2][14][15]<=-140; ws[2][14][16]<=-109; ws[2][14][17]<= -65; ws[2][14][18]<=  61; ws[2][14][19]<= 124; ws[2][14][20]<=  75; ws[2][14][21]<= -71; ws[2][14][22]<=-105; ws[2][14][23]<= -49; ws[2][14][24]<=  22; ws[2][14][25]<= 172; ws[2][14][26]<= 186; ws[2][14][27]<=  43; ws[2][14][28]<=   9; ws[2][14][29]<= -87; ws[2][14][30]<=  27; ws[2][14][31]<= 159; ws[2][14][32]<= 243; ws[2][14][33]<= 208; ws[2][14][34]<=  36; ws[2][14][35]<= -15; ws[2][14][36]<=  69; ws[2][14][37]<=  57; ws[2][14][38]<= 149; ws[2][14][39]<= 203; ws[2][14][40]<= 172; ws[2][14][41]<=   7; ws[2][14][42]<=  27; ws[2][14][43]<=  42; ws[2][14][44]<=  51; ws[2][14][45]<= 175; ws[2][14][46]<= 211; ws[2][14][47]<= 184; ws[2][14][48]<=  78;
        ws[2][15][0]<=  63; ws[2][15][1]<=  79; ws[2][15][2]<=  52; ws[2][15][3]<= -61; ws[2][15][4]<= -68; ws[2][15][5]<= -25; ws[2][15][6]<=  45; ws[2][15][7]<=  84; ws[2][15][8]<= 106; ws[2][15][9]<=-113; ws[2][15][10]<=-152; ws[2][15][11]<= -47; ws[2][15][12]<=  42; ws[2][15][13]<= 135; ws[2][15][14]<=  93; ws[2][15][15]<=   5; ws[2][15][16]<=-143; ws[2][15][17]<= -64; ws[2][15][18]<= 120; ws[2][15][19]<= 198; ws[2][15][20]<= 130; ws[2][15][21]<=  54; ws[2][15][22]<=   2; ws[2][15][23]<=-116; ws[2][15][24]<= -10; ws[2][15][25]<= 150; ws[2][15][26]<= 179; ws[2][15][27]<=  43; ws[2][15][28]<=  68; ws[2][15][29]<= -29; ws[2][15][30]<=   4; ws[2][15][31]<= 115; ws[2][15][32]<= 190; ws[2][15][33]<= 188; ws[2][15][34]<=  25; ws[2][15][35]<=   6; ws[2][15][36]<= -16; ws[2][15][37]<=  13; ws[2][15][38]<= 116; ws[2][15][39]<= 140; ws[2][15][40]<=  88; ws[2][15][41]<= -53; ws[2][15][42]<= -77; ws[2][15][43]<= -73; ws[2][15][44]<=  11; ws[2][15][45]<=  21; ws[2][15][46]<= 108; ws[2][15][47]<=  19; ws[2][15][48]<=  37;

        ws[3][0 ][0]<=-113; ws[3][0 ][1]<= 175; ws[3][0 ][2]<= 181; ws[3][0 ][3]<= 127; ws[3][0 ][4]<= -19; ws[3][0 ][5]<=-140; ws[3][0 ][6]<=-246; ws[3][0 ][7]<= -73; ws[3][0 ][8]<=  76; ws[3][0 ][9]<= 136; ws[3][0 ][10]<= 102; ws[3][0 ][11]<= -73; ws[3][0 ][12]<= -93; ws[3][0 ][13]<=-212; ws[3][0 ][14]<= -74; ws[3][0 ][15]<=  42; ws[3][0 ][16]<=  53; ws[3][0 ][17]<=  84; ws[3][0 ][18]<= -65; ws[3][0 ][19]<= -91; ws[3][0 ][20]<= -97; ws[3][0 ][21]<=-108; ws[3][0 ][22]<= -99; ws[3][0 ][23]<=  29; ws[3][0 ][24]<=  94; ws[3][0 ][25]<= -47; ws[3][0 ][26]<= -23; ws[3][0 ][27]<= -45; ws[3][0 ][28]<= -57; ws[3][0 ][29]<=-122; ws[3][0 ][30]<=  60; ws[3][0 ][31]<= 103; ws[3][0 ][32]<= -20; ws[3][0 ][33]<= -46; ws[3][0 ][34]<= -24; ws[3][0 ][35]<=  83; ws[3][0 ][36]<= -70; ws[3][0 ][37]<=   3; ws[3][0 ][38]<=  54; ws[3][0 ][39]<=  -5; ws[3][0 ][40]<=-131; ws[3][0 ][41]<= -32; ws[3][0 ][42]<= 205; ws[3][0 ][43]<=  57; ws[3][0 ][44]<=  55; ws[3][0 ][45]<=  55; ws[3][0 ][46]<= -41; ws[3][0 ][47]<=-131; ws[3][0 ][48]<=-119;
        ws[3][1 ][0]<=  23; ws[3][1 ][1]<=  39; ws[3][1 ][2]<=  36; ws[3][1 ][3]<=  92; ws[3][1 ][4]<=   4; ws[3][1 ][5]<=  -1; ws[3][1 ][6]<=  73; ws[3][1 ][7]<=  67; ws[3][1 ][8]<=   1; ws[3][1 ][9]<=  79; ws[3][1 ][10]<=  95; ws[3][1 ][11]<=  57; ws[3][1 ][12]<=  59; ws[3][1 ][13]<=  79; ws[3][1 ][14]<=  31; ws[3][1 ][15]<=  77; ws[3][1 ][16]<=  39; ws[3][1 ][17]<=  71; ws[3][1 ][18]<=  36; ws[3][1 ][19]<=  79; ws[3][1 ][20]<=  34; ws[3][1 ][21]<=  91; ws[3][1 ][22]<=  87; ws[3][1 ][23]<=  94; ws[3][1 ][24]<=  42; ws[3][1 ][25]<=  13; ws[3][1 ][26]<=  20; ws[3][1 ][27]<=  60; ws[3][1 ][28]<=  61; ws[3][1 ][29]<=  85; ws[3][1 ][30]<=  52; ws[3][1 ][31]<=  46; ws[3][1 ][32]<=  31; ws[3][1 ][33]<=  92; ws[3][1 ][34]<=  31; ws[3][1 ][35]<=  99; ws[3][1 ][36]<=  91; ws[3][1 ][37]<=  27; ws[3][1 ][38]<=  53; ws[3][1 ][39]<=  80; ws[3][1 ][40]<=  70; ws[3][1 ][41]<=  47; ws[3][1 ][42]<=  68; ws[3][1 ][43]<=  30; ws[3][1 ][44]<=  97; ws[3][1 ][45]<=  57; ws[3][1 ][46]<=  94; ws[3][1 ][47]<=  14; ws[3][1 ][48]<=  45;
        ws[3][2 ][0]<= -16; ws[3][2 ][1]<=   9; ws[3][2 ][2]<=  18; ws[3][2 ][3]<=  55; ws[3][2 ][4]<= -24; ws[3][2 ][5]<=   2; ws[3][2 ][6]<= -40; ws[3][2 ][7]<=  12; ws[3][2 ][8]<=  39; ws[3][2 ][9]<= 109; ws[3][2 ][10]<= 129; ws[3][2 ][11]<=  71; ws[3][2 ][12]<=  19; ws[3][2 ][13]<= -55; ws[3][2 ][14]<=  49; ws[3][2 ][15]<=  84; ws[3][2 ][16]<= 154; ws[3][2 ][17]<= 176; ws[3][2 ][18]<= 103; ws[3][2 ][19]<=  -8; ws[3][2 ][20]<= -70; ws[3][2 ][21]<=  62; ws[3][2 ][22]<= 110; ws[3][2 ][23]<= 171; ws[3][2 ][24]<= 206; ws[3][2 ][25]<= 114; ws[3][2 ][26]<=  63; ws[3][2 ][27]<=   3; ws[3][2 ][28]<=  26; ws[3][2 ][29]<=  88; ws[3][2 ][30]<= 114; ws[3][2 ][31]<= 174; ws[3][2 ][32]<=  93; ws[3][2 ][33]<=  62; ws[3][2 ][34]<= -82; ws[3][2 ][35]<=  44; ws[3][2 ][36]<=  -8; ws[3][2 ][37]<= 120; ws[3][2 ][38]<= 111; ws[3][2 ][39]<=  85; ws[3][2 ][40]<= -15; ws[3][2 ][41]<= -79; ws[3][2 ][42]<= -67; ws[3][2 ][43]<= -54; ws[3][2 ][44]<=  -7; ws[3][2 ][45]<=  53; ws[3][2 ][46]<=  23; ws[3][2 ][47]<= -12; ws[3][2 ][48]<=-135;
        ws[3][3 ][0]<= -57; ws[3][3 ][1]<=  74; ws[3][3 ][2]<= 184; ws[3][3 ][3]<=  74; ws[3][3 ][4]<=-104; ws[3][3 ][5]<= -18; ws[3][3 ][6]<=  83; ws[3][3 ][7]<=-106; ws[3][3 ][8]<=  27; ws[3][3 ][9]<= 108; ws[3][3 ][10]<=  49; ws[3][3 ][11]<= -12; ws[3][3 ][12]<=  22; ws[3][3 ][13]<= 124; ws[3][3 ][14]<=-168; ws[3][3 ][15]<= -73; ws[3][3 ][16]<=  27; ws[3][3 ][17]<= 134; ws[3][3 ][18]<=  27; ws[3][3 ][19]<= 103; ws[3][3 ][20]<= 119; ws[3][3 ][21]<=-195; ws[3][3 ][22]<=-175; ws[3][3 ][23]<= -43; ws[3][3 ][24]<= 122; ws[3][3 ][25]<= 147; ws[3][3 ][26]<= 112; ws[3][3 ][27]<=  92; ws[3][3 ][28]<=-132; ws[3][3 ][29]<=-226; ws[3][3 ][30]<=-111; ws[3][3 ][31]<= 110; ws[3][3 ][32]<= 134; ws[3][3 ][33]<= 131; ws[3][3 ][34]<=  97; ws[3][3 ][35]<= -19; ws[3][3 ][36]<=-168; ws[3][3 ][37]<=-111; ws[3][3 ][38]<=  54; ws[3][3 ][39]<= 122; ws[3][3 ][40]<=  85; ws[3][3 ][41]<=  38; ws[3][3 ][42]<=  31; ws[3][3 ][43]<= -39; ws[3][3 ][44]<=-171; ws[3][3 ][45]<= -57; ws[3][3 ][46]<= 114; ws[3][3 ][47]<=  26; ws[3][3 ][48]<=  77;
        ws[3][4 ][0]<=  19; ws[3][4 ][1]<=  82; ws[3][4 ][2]<=  41; ws[3][4 ][3]<= -76; ws[3][4 ][4]<=-157; ws[3][4 ][5]<=-106; ws[3][4 ][6]<=-106; ws[3][4 ][7]<=  90; ws[3][4 ][8]<=  88; ws[3][4 ][9]<=   4; ws[3][4 ][10]<=-104; ws[3][4 ][11]<=-213; ws[3][4 ][12]<=-149; ws[3][4 ][13]<=-108; ws[3][4 ][14]<= 103; ws[3][4 ][15]<= 107; ws[3][4 ][16]<=  46; ws[3][4 ][17]<= -15; ws[3][4 ][18]<=-155; ws[3][4 ][19]<=-140; ws[3][4 ][20]<=-168; ws[3][4 ][21]<= 119; ws[3][4 ][22]<=  85; ws[3][4 ][23]<=  97; ws[3][4 ][24]<= -11; ws[3][4 ][25]<= -89; ws[3][4 ][26]<=-159; ws[3][4 ][27]<=-122; ws[3][4 ][28]<=  53; ws[3][4 ][29]<=  23; ws[3][4 ][30]<= 138; ws[3][4 ][31]<= 110; ws[3][4 ][32]<= -23; ws[3][4 ][33]<= -43; ws[3][4 ][34]<= -94; ws[3][4 ][35]<=  87; ws[3][4 ][36]<= -10; ws[3][4 ][37]<=  61; ws[3][4 ][38]<= 157; ws[3][4 ][39]<=  87; ws[3][4 ][40]<= -45; ws[3][4 ][41]<=  -7; ws[3][4 ][42]<=  19; ws[3][4 ][43]<= -60; ws[3][4 ][44]<=  32; ws[3][4 ][45]<=  76; ws[3][4 ][46]<=  63; ws[3][4 ][47]<=  10; ws[3][4 ][48]<= -54;
        ws[3][5 ][0]<= -87; ws[3][5 ][1]<=  38; ws[3][5 ][2]<= 155; ws[3][5 ][3]<=  70; ws[3][5 ][4]<= -18; ws[3][5 ][5]<=-171; ws[3][5 ][6]<=-196; ws[3][5 ][7]<= -82; ws[3][5 ][8]<=  42; ws[3][5 ][9]<= 141; ws[3][5 ][10]<= 105; ws[3][5 ][11]<= -72; ws[3][5 ][12]<=-175; ws[3][5 ][13]<=-147; ws[3][5 ][14]<= -29; ws[3][5 ][15]<=  97; ws[3][5 ][16]<= 113; ws[3][5 ][17]<=  83; ws[3][5 ][18]<= -87; ws[3][5 ][19]<=-102; ws[3][5 ][20]<=-113; ws[3][5 ][21]<= -56; ws[3][5 ][22]<=  58; ws[3][5 ][23]<= 129; ws[3][5 ][24]<=  73; ws[3][5 ][25]<=-107; ws[3][5 ][26]<= -80; ws[3][5 ][27]<= -98; ws[3][5 ][28]<=  -8; ws[3][5 ][29]<=  36; ws[3][5 ][30]<=  75; ws[3][5 ][31]<=  -1; ws[3][5 ][32]<=-110; ws[3][5 ][33]<=-150; ws[3][5 ][34]<= -83; ws[3][5 ][35]<= -59; ws[3][5 ][36]<=  18; ws[3][5 ][37]<=  79; ws[3][5 ][38]<=  -7; ws[3][5 ][39]<= -93; ws[3][5 ][40]<=-168; ws[3][5 ][41]<=-113; ws[3][5 ][42]<= -43; ws[3][5 ][43]<=  34; ws[3][5 ][44]<=  68; ws[3][5 ][45]<= -52; ws[3][5 ][46]<=-185; ws[3][5 ][47]<=-190; ws[3][5 ][48]<= -75;
        ws[3][6 ][0]<=  57; ws[3][6 ][1]<=  -6; ws[3][6 ][2]<= -17; ws[3][6 ][3]<=  98; ws[3][6 ][4]<=  21; ws[3][6 ][5]<=   6; ws[3][6 ][6]<=  38; ws[3][6 ][7]<=  38; ws[3][6 ][8]<=  -8; ws[3][6 ][9]<=  16; ws[3][6 ][10]<= 108; ws[3][6 ][11]<=  70; ws[3][6 ][12]<=  47; ws[3][6 ][13]<=   0; ws[3][6 ][14]<=  31; ws[3][6 ][15]<=  -2; ws[3][6 ][16]<=  49; ws[3][6 ][17]<= 140; ws[3][6 ][18]<=  75; ws[3][6 ][19]<=  46; ws[3][6 ][20]<=  50; ws[3][6 ][21]<=  59; ws[3][6 ][22]<= -24; ws[3][6 ][23]<=  64; ws[3][6 ][24]<= 162; ws[3][6 ][25]<= 121; ws[3][6 ][26]<=  41; ws[3][6 ][27]<=  91; ws[3][6 ][28]<=  28; ws[3][6 ][29]<=  72; ws[3][6 ][30]<=  68; ws[3][6 ][31]<= 163; ws[3][6 ][32]<= 106; ws[3][6 ][33]<=  22; ws[3][6 ][34]<=  61; ws[3][6 ][35]<=  78; ws[3][6 ][36]<=  75; ws[3][6 ][37]<=  95; ws[3][6 ][38]<= 214; ws[3][6 ][39]<= 152; ws[3][6 ][40]<=  53; ws[3][6 ][41]<=  16; ws[3][6 ][42]<= 190; ws[3][6 ][43]<= 116; ws[3][6 ][44]<= 152; ws[3][6 ][45]<= 237; ws[3][6 ][46]<= 135; ws[3][6 ][47]<=  82; ws[3][6 ][48]<=  83;
        ws[3][7 ][0]<= -30; ws[3][7 ][1]<= -84; ws[3][7 ][2]<=-167; ws[3][7 ][3]<=-148; ws[3][7 ][4]<= -95; ws[3][7 ][5]<=  26; ws[3][7 ][6]<= 129; ws[3][7 ][7]<= 121; ws[3][7 ][8]<= -72; ws[3][7 ][9]<=-103; ws[3][7 ][10]<=-131; ws[3][7 ][11]<= -75; ws[3][7 ][12]<= -36; ws[3][7 ][13]<= 107; ws[3][7 ][14]<= 150; ws[3][7 ][15]<=  34; ws[3][7 ][16]<= -61; ws[3][7 ][17]<=-109; ws[3][7 ][18]<= -43; ws[3][7 ][19]<= -25; ws[3][7 ][20]<=  94; ws[3][7 ][21]<= 191; ws[3][7 ][22]<=  96; ws[3][7 ][23]<= -16; ws[3][7 ][24]<= -99; ws[3][7 ][25]<= -32; ws[3][7 ][26]<=  24; ws[3][7 ][27]<= 102; ws[3][7 ][28]<= 232; ws[3][7 ][29]<= 186; ws[3][7 ][30]<=  29; ws[3][7 ][31]<= -79; ws[3][7 ][32]<=  -3; ws[3][7 ][33]<=  29; ws[3][7 ][34]<=  55; ws[3][7 ][35]<= 152; ws[3][7 ][36]<= 129; ws[3][7 ][37]<= 101; ws[3][7 ][38]<=  30; ws[3][7 ][39]<=  -8; ws[3][7 ][40]<=  76; ws[3][7 ][41]<=  72; ws[3][7 ][42]<= -33; ws[3][7 ][43]<=  19; ws[3][7 ][44]<=  91; ws[3][7 ][45]<=  22; ws[3][7 ][46]<= -30; ws[3][7 ][47]<=  52; ws[3][7 ][48]<= 121;
        ws[3][8 ][0]<=-204; ws[3][8 ][1]<=-145; ws[3][8 ][2]<= -99; ws[3][8 ][3]<=-138; ws[3][8 ][4]<=-135; ws[3][8 ][5]<= -81; ws[3][8 ][6]<=-146; ws[3][8 ][7]<=-129; ws[3][8 ][8]<= -81; ws[3][8 ][9]<= -59; ws[3][8 ][10]<= -41; ws[3][8 ][11]<=-105; ws[3][8 ][12]<=-119; ws[3][8 ][13]<=-145; ws[3][8 ][14]<= -31; ws[3][8 ][15]<=-108; ws[3][8 ][16]<= -63; ws[3][8 ][17]<=   3; ws[3][8 ][18]<= -45; ws[3][8 ][19]<=-101; ws[3][8 ][20]<=-114; ws[3][8 ][21]<= -61; ws[3][8 ][22]<=-113; ws[3][8 ][23]<=  38; ws[3][8 ][24]<=  27; ws[3][8 ][25]<= -68; ws[3][8 ][26]<= -63; ws[3][8 ][27]<= -28; ws[3][8 ][28]<= -93; ws[3][8 ][29]<=-116; ws[3][8 ][30]<=  21; ws[3][8 ][31]<=  54; ws[3][8 ][32]<=   9; ws[3][8 ][33]<= -14; ws[3][8 ][34]<=   3; ws[3][8 ][35]<= -41; ws[3][8 ][36]<= -95; ws[3][8 ][37]<=   0; ws[3][8 ][38]<=  15; ws[3][8 ][39]<=  -8; ws[3][8 ][40]<= -33; ws[3][8 ][41]<=  12; ws[3][8 ][42]<= -47; ws[3][8 ][43]<=-177; ws[3][8 ][44]<=-144; ws[3][8 ][45]<= -19; ws[3][8 ][46]<=  23; ws[3][8 ][47]<= -25; ws[3][8 ][48]<=  -8;
        ws[3][9 ][0]<=  30; ws[3][9 ][1]<= -99; ws[3][9 ][2]<=-200; ws[3][9 ][3]<=-181; ws[3][9 ][4]<=-146; ws[3][9 ][5]<= -32; ws[3][9 ][6]<= -29; ws[3][9 ][7]<=  -7; ws[3][9 ][8]<=  16; ws[3][9 ][9]<= -10; ws[3][9 ][10]<= -45; ws[3][9 ][11]<= -59; ws[3][9 ][12]<= -55; ws[3][9 ][13]<=   0; ws[3][9 ][14]<=  33; ws[3][9 ][15]<= 107; ws[3][9 ][16]<= 119; ws[3][9 ][17]<=  51; ws[3][9 ][18]<= -63; ws[3][9 ][19]<=-106; ws[3][9 ][20]<= -48; ws[3][9 ][21]<=  66; ws[3][9 ][22]<= 150; ws[3][9 ][23]<= 105; ws[3][9 ][24]<= -47; ws[3][9 ][25]<=-127; ws[3][9 ][26]<= -54; ws[3][9 ][27]<=   5; ws[3][9 ][28]<=  70; ws[3][9 ][29]<=  93; ws[3][9 ][30]<=  57; ws[3][9 ][31]<=-119; ws[3][9 ][32]<= -85; ws[3][9 ][33]<= -38; ws[3][9 ][34]<= 146; ws[3][9 ][35]<=  23; ws[3][9 ][36]<=  53; ws[3][9 ][37]<= -88; ws[3][9 ][38]<=-125; ws[3][9 ][39]<= -63; ws[3][9 ][40]<= 149; ws[3][9 ][41]<= 226; ws[3][9 ][42]<=  10; ws[3][9 ][43]<= -69; ws[3][9 ][44]<=-147; ws[3][9 ][45]<=-188; ws[3][9 ][46]<= -10; ws[3][9 ][47]<= 226; ws[3][9 ][48]<= 244;
        ws[3][10][0]<=  52; ws[3][10][1]<= -27; ws[3][10][2]<= -88; ws[3][10][3]<= -48; ws[3][10][4]<=-108; ws[3][10][5]<=-111; ws[3][10][6]<=-188; ws[3][10][7]<= 125; ws[3][10][8]<= -17; ws[3][10][9]<= -58; ws[3][10][10]<= -84; ws[3][10][11]<=-122; ws[3][10][12]<=-134; ws[3][10][13]<=-130; ws[3][10][14]<=  42; ws[3][10][15]<= -16; ws[3][10][16]<= -22; ws[3][10][17]<= -93; ws[3][10][18]<= -66; ws[3][10][19]<=-137; ws[3][10][20]<=-178; ws[3][10][21]<=  46; ws[3][10][22]<= -50; ws[3][10][23]<= -72; ws[3][10][24]<= -18; ws[3][10][25]<= -69; ws[3][10][26]<=-136; ws[3][10][27]<= -70; ws[3][10][28]<=-103; ws[3][10][29]<= -88; ws[3][10][30]<= -57; ws[3][10][31]<= -84; ws[3][10][32]<= -72; ws[3][10][33]<= -75; ws[3][10][34]<=-102; ws[3][10][35]<=-167; ws[3][10][36]<=-150; ws[3][10][37]<= -52; ws[3][10][38]<= -54; ws[3][10][39]<=  -8; ws[3][10][40]<= -76; ws[3][10][41]<=-123; ws[3][10][42]<=-263; ws[3][10][43]<=-162; ws[3][10][44]<= -35; ws[3][10][45]<= -74; ws[3][10][46]<= -15; ws[3][10][47]<= -29; ws[3][10][48]<=-135;
        ws[3][11][0]<= -37; ws[3][11][1]<=-127; ws[3][11][2]<=-149; ws[3][11][3]<= -46; ws[3][11][4]<= -14; ws[3][11][5]<=  31; ws[3][11][6]<=  31; ws[3][11][7]<=  32; ws[3][11][8]<= -94; ws[3][11][9]<=-149; ws[3][11][10]<= -31; ws[3][11][11]<=  -9; ws[3][11][12]<=  26; ws[3][11][13]<=  35; ws[3][11][14]<=  64; ws[3][11][15]<= -43; ws[3][11][16]<=-165; ws[3][11][17]<= -64; ws[3][11][18]<= -10; ws[3][11][19]<=   3; ws[3][11][20]<=  40; ws[3][11][21]<= -14; ws[3][11][22]<=-117; ws[3][11][23]<= -73; ws[3][11][24]<= -75; ws[3][11][25]<= -27; ws[3][11][26]<=  10; ws[3][11][27]<= -28; ws[3][11][28]<=   1; ws[3][11][29]<= -96; ws[3][11][30]<=-142; ws[3][11][31]<= -58; ws[3][11][32]<= -11; ws[3][11][33]<=  33; ws[3][11][34]<=  29; ws[3][11][35]<= -89; ws[3][11][36]<=-129; ws[3][11][37]<=-120; ws[3][11][38]<=   8; ws[3][11][39]<=  31; ws[3][11][40]<=  19; ws[3][11][41]<=  -1; ws[3][11][42]<=-163; ws[3][11][43]<=-108; ws[3][11][44]<= -63; ws[3][11][45]<=  50; ws[3][11][46]<=  42; ws[3][11][47]<=  69; ws[3][11][48]<=  30;
        ws[3][12][0]<=  84; ws[3][12][1]<=  67; ws[3][12][2]<= -47; ws[3][12][3]<=-152; ws[3][12][4]<=-147; ws[3][12][5]<= -97; ws[3][12][6]<=-113; ws[3][12][7]<=  68; ws[3][12][8]<= 128; ws[3][12][9]<=  76; ws[3][12][10]<= -97; ws[3][12][11]<=-167; ws[3][12][12]<=-159; ws[3][12][13]<=-136; ws[3][12][14]<= -15; ws[3][12][15]<=  70; ws[3][12][16]<=  96; ws[3][12][17]<= -15; ws[3][12][18]<=-140; ws[3][12][19]<=-117; ws[3][12][20]<=-133; ws[3][12][21]<= -48; ws[3][12][22]<=  54; ws[3][12][23]<=  67; ws[3][12][24]<= 108; ws[3][12][25]<= -54; ws[3][12][26]<= -99; ws[3][12][27]<=-116; ws[3][12][28]<= -41; ws[3][12][29]<= -53; ws[3][12][30]<=  42; ws[3][12][31]<= 150; ws[3][12][32]<= 130; ws[3][12][33]<=  11; ws[3][12][34]<= -45; ws[3][12][35]<= -30; ws[3][12][36]<= -60; ws[3][12][37]<=  51; ws[3][12][38]<= 250; ws[3][12][39]<= 237; ws[3][12][40]<=  64; ws[3][12][41]<=   3; ws[3][12][42]<=  81; ws[3][12][43]<= -58; ws[3][12][44]<=  41; ws[3][12][45]<= 215; ws[3][12][46]<= 286; ws[3][12][47]<= 140; ws[3][12][48]<= -57;
        ws[3][13][0]<= 201; ws[3][13][1]<= 175; ws[3][13][2]<=  41; ws[3][13][3]<= -59; ws[3][13][4]<=-139; ws[3][13][5]<= -64; ws[3][13][6]<= -82; ws[3][13][7]<=  98; ws[3][13][8]<= 168; ws[3][13][9]<=  70; ws[3][13][10]<= -25; ws[3][13][11]<=-126; ws[3][13][12]<=-146; ws[3][13][13]<=-108; ws[3][13][14]<=  98; ws[3][13][15]<= 129; ws[3][13][16]<=  71; ws[3][13][17]<=-103; ws[3][13][18]<= -70; ws[3][13][19]<=-132; ws[3][13][20]<= -70; ws[3][13][21]<=  18; ws[3][13][22]<=  84; ws[3][13][23]<=  58; ws[3][13][24]<= -41; ws[3][13][25]<=-117; ws[3][13][26]<=-120; ws[3][13][27]<= -82; ws[3][13][28]<=  55; ws[3][13][29]<=  90; ws[3][13][30]<=  24; ws[3][13][31]<=  18; ws[3][13][32]<= -31; ws[3][13][33]<=  -1; ws[3][13][34]<= -22; ws[3][13][35]<=  90; ws[3][13][36]<=  66; ws[3][13][37]<=   7; ws[3][13][38]<= -26; ws[3][13][39]<= -35; ws[3][13][40]<=  27; ws[3][13][41]<= -27; ws[3][13][42]<= 122; ws[3][13][43]<=  87; ws[3][13][44]<=  93; ws[3][13][45]<=   0; ws[3][13][46]<=  43; ws[3][13][47]<=  -9; ws[3][13][48]<=  64;
        ws[3][14][0]<=  80; ws[3][14][1]<=  -2; ws[3][14][2]<= -60; ws[3][14][3]<=-125; ws[3][14][4]<= -74; ws[3][14][5]<= -74; ws[3][14][6]<=  50; ws[3][14][7]<=  50; ws[3][14][8]<= -52; ws[3][14][9]<= -68; ws[3][14][10]<=-169; ws[3][14][11]<=-158; ws[3][14][12]<= -71; ws[3][14][13]<=  19; ws[3][14][14]<=  -9; ws[3][14][15]<=  15; ws[3][14][16]<= -69; ws[3][14][17]<=-110; ws[3][14][18]<=-167; ws[3][14][19]<=-128; ws[3][14][20]<= -24; ws[3][14][21]<=  19; ws[3][14][22]<=  55; ws[3][14][23]<=  -3; ws[3][14][24]<= -68; ws[3][14][25]<= -81; ws[3][14][26]<= -89; ws[3][14][27]<=  15; ws[3][14][28]<=  99; ws[3][14][29]<=  66; ws[3][14][30]<=  -9; ws[3][14][31]<=-105; ws[3][14][32]<= -79; ws[3][14][33]<= -77; ws[3][14][34]<= -19; ws[3][14][35]<= 126; ws[3][14][36]<= 102; ws[3][14][37]<= -10; ws[3][14][38]<= -74; ws[3][14][39]<= -69; ws[3][14][40]<= -77; ws[3][14][41]<=   7; ws[3][14][42]<= 186; ws[3][14][43]<= 176; ws[3][14][44]<=  26; ws[3][14][45]<= -70; ws[3][14][46]<=-121; ws[3][14][47]<=-125; ws[3][14][48]<= -22;
        ws[3][15][0]<=  50; ws[3][15][1]<=  35; ws[3][15][2]<=  62; ws[3][15][3]<=  50; ws[3][15][4]<=  81; ws[3][15][5]<= -11; ws[3][15][6]<= -59; ws[3][15][7]<=  15; ws[3][15][8]<= -72; ws[3][15][9]<=  -7; ws[3][15][10]<= 126; ws[3][15][11]<= 141; ws[3][15][12]<=  48; ws[3][15][13]<= -50; ws[3][15][14]<=  40; ws[3][15][15]<=  14; ws[3][15][16]<=  42; ws[3][15][17]<=  94; ws[3][15][18]<= 137; ws[3][15][19]<=  27; ws[3][15][20]<= -14; ws[3][15][21]<=  32; ws[3][15][22]<=  -7; ws[3][15][23]<=  79; ws[3][15][24]<=  66; ws[3][15][25]<=  61; ws[3][15][26]<= -78; ws[3][15][27]<=-117; ws[3][15][28]<= 116; ws[3][15][29]<=   3; ws[3][15][30]<= -55; ws[3][15][31]<= -96; ws[3][15][32]<=-172; ws[3][15][33]<=-113; ws[3][15][34]<=-115; ws[3][15][35]<= 102; ws[3][15][36]<= -22; ws[3][15][37]<= -99; ws[3][15][38]<=-210; ws[3][15][39]<=-206; ws[3][15][40]<=-146; ws[3][15][41]<= -50; ws[3][15][42]<= 121; ws[3][15][43]<= -37; ws[3][15][44]<=-144; ws[3][15][45]<=-228; ws[3][15][46]<=-217; ws[3][15][47]<=-118; ws[3][15][48]<= -85;

        ws[4][0 ][0]<= 157; ws[4][0 ][1]<=  83; ws[4][0 ][2]<=  74; ws[4][0 ][3]<= 221; ws[4][0 ][4]<=  63; ws[4][0 ][5]<= -44; ws[4][0 ][6]<= -34; ws[4][0 ][7]<= 156; ws[4][0 ][8]<= 105; ws[4][0 ][9]<=  81; ws[4][0 ][10]<= 111; ws[4][0 ][11]<=  71; ws[4][0 ][12]<=-156; ws[4][0 ][13]<=-151; ws[4][0 ][14]<=  93; ws[4][0 ][15]<=  53; ws[4][0 ][16]<=  27; ws[4][0 ][17]<= 111; ws[4][0 ][18]<=  83; ws[4][0 ][19]<=-141; ws[4][0 ][20]<=-224; ws[4][0 ][21]<=  38; ws[4][0 ][22]<=  -5; ws[4][0 ][23]<= -80; ws[4][0 ][24]<=  48; ws[4][0 ][25]<= 102; ws[4][0 ][26]<= -76; ws[4][0 ][27]<=-179; ws[4][0 ][28]<=  27; ws[4][0 ][29]<= -80; ws[4][0 ][30]<= -61; ws[4][0 ][31]<=  15; ws[4][0 ][32]<= 100; ws[4][0 ][33]<= -48; ws[4][0 ][34]<=-165; ws[4][0 ][35]<=  -1; ws[4][0 ][36]<= -59; ws[4][0 ][37]<=-110; ws[4][0 ][38]<=-105; ws[4][0 ][39]<=  62; ws[4][0 ][40]<=  86; ws[4][0 ][41]<=  -5; ws[4][0 ][42]<= -71; ws[4][0 ][43]<= -42; ws[4][0 ][44]<= -85; ws[4][0 ][45]<=-101; ws[4][0 ][46]<=   8; ws[4][0 ][47]<=  90; ws[4][0 ][48]<=  41;
        ws[4][1 ][0]<=-112; ws[4][1 ][1]<=  32; ws[4][1 ][2]<=  15; ws[4][1 ][3]<= -41; ws[4][1 ][4]<= -28; ws[4][1 ][5]<=  80; ws[4][1 ][6]<= 142; ws[4][1 ][7]<= -46; ws[4][1 ][8]<= -16; ws[4][1 ][9]<= -11; ws[4][1 ][10]<= -27; ws[4][1 ][11]<=  43; ws[4][1 ][12]<=  70; ws[4][1 ][13]<= 258; ws[4][1 ][14]<= -18; ws[4][1 ][15]<=  54; ws[4][1 ][16]<=  52; ws[4][1 ][17]<=  46; ws[4][1 ][18]<=  85; ws[4][1 ][19]<=  75; ws[4][1 ][20]<= 210; ws[4][1 ][21]<=  26; ws[4][1 ][22]<=  51; ws[4][1 ][23]<=  57; ws[4][1 ][24]<=  37; ws[4][1 ][25]<=  86; ws[4][1 ][26]<= 142; ws[4][1 ][27]<= 250; ws[4][1 ][28]<=  17; ws[4][1 ][29]<= 122; ws[4][1 ][30]<=  65; ws[4][1 ][31]<=  49; ws[4][1 ][32]<=  46; ws[4][1 ][33]<= 121; ws[4][1 ][34]<= 280; ws[4][1 ][35]<=   4; ws[4][1 ][36]<=  90; ws[4][1 ][37]<=  97; ws[4][1 ][38]<=  82; ws[4][1 ][39]<=  54; ws[4][1 ][40]<= 147; ws[4][1 ][41]<= 301; ws[4][1 ][42]<=  18; ws[4][1 ][43]<= 127; ws[4][1 ][44]<=  97; ws[4][1 ][45]<=  71; ws[4][1 ][46]<=  58; ws[4][1 ][47]<= 158; ws[4][1 ][48]<= 271;
        ws[4][2 ][0]<= -31; ws[4][2 ][1]<= -30; ws[4][2 ][2]<= -16; ws[4][2 ][3]<= -23; ws[4][2 ][4]<=-160; ws[4][2 ][5]<=-259; ws[4][2 ][6]<=-146; ws[4][2 ][7]<= -25; ws[4][2 ][8]<=  -9; ws[4][2 ][9]<=  75; ws[4][2 ][10]<= -23; ws[4][2 ][11]<=-206; ws[4][2 ][12]<=-205; ws[4][2 ][13]<=-123; ws[4][2 ][14]<=  21; ws[4][2 ][15]<=  17; ws[4][2 ][16]<=  46; ws[4][2 ][17]<= -94; ws[4][2 ][18]<=-116; ws[4][2 ][19]<= -99; ws[4][2 ][20]<=-109; ws[4][2 ][21]<= -37; ws[4][2 ][22]<= -28; ws[4][2 ][23]<= -87; ws[4][2 ][24]<= -60; ws[4][2 ][25]<= -79; ws[4][2 ][26]<= -13; ws[4][2 ][27]<=  65; ws[4][2 ][28]<= -44; ws[4][2 ][29]<= -60; ws[4][2 ][30]<= -53; ws[4][2 ][31]<=  11; ws[4][2 ][32]<= 112; ws[4][2 ][33]<= 110; ws[4][2 ][34]<=  89; ws[4][2 ][35]<= -29; ws[4][2 ][36]<=-105; ws[4][2 ][37]<=  -3; ws[4][2 ][38]<= 117; ws[4][2 ][39]<= 180; ws[4][2 ][40]<= 211; ws[4][2 ][41]<= 182; ws[4][2 ][42]<=  52; ws[4][2 ][43]<=  11; ws[4][2 ][44]<=  98; ws[4][2 ][45]<= 255; ws[4][2 ][46]<= 276; ws[4][2 ][47]<= 212; ws[4][2 ][48]<= 145;
        ws[4][3 ][0]<=-119; ws[4][3 ][1]<= -78; ws[4][3 ][2]<= -89; ws[4][3 ][3]<=  40; ws[4][3 ][4]<= 115; ws[4][3 ][5]<= 115; ws[4][3 ][6]<= 105; ws[4][3 ][7]<= -78; ws[4][3 ][8]<= -43; ws[4][3 ][9]<= -11; ws[4][3 ][10]<=   4; ws[4][3 ][11]<=  72; ws[4][3 ][12]<= 114; ws[4][3 ][13]<=  78; ws[4][3 ][14]<=-118; ws[4][3 ][15]<= -52; ws[4][3 ][16]<= -69; ws[4][3 ][17]<=   0; ws[4][3 ][18]<=  86; ws[4][3 ][19]<= 125; ws[4][3 ][20]<=  44; ws[4][3 ][21]<= -45; ws[4][3 ][22]<= -30; ws[4][3 ][23]<=  19; ws[4][3 ][24]<=  78; ws[4][3 ][25]<=  50; ws[4][3 ][26]<= 122; ws[4][3 ][27]<=  36; ws[4][3 ][28]<= -64; ws[4][3 ][29]<= -33; ws[4][3 ][30]<=  50; ws[4][3 ][31]<=  39; ws[4][3 ][32]<= 129; ws[4][3 ][33]<=  91; ws[4][3 ][34]<=   6; ws[4][3 ][35]<=-113; ws[4][3 ][36]<=  -2; ws[4][3 ][37]<=  53; ws[4][3 ][38]<= 112; ws[4][3 ][39]<= 123; ws[4][3 ][40]<=  94; ws[4][3 ][41]<=  12; ws[4][3 ][42]<=-116; ws[4][3 ][43]<= -10; ws[4][3 ][44]<=  97; ws[4][3 ][45]<= 103; ws[4][3 ][46]<=  62; ws[4][3 ][47]<=  82; ws[4][3 ][48]<=  43;
        ws[4][4 ][0]<=   2; ws[4][4 ][1]<=  70; ws[4][4 ][2]<= 114; ws[4][4 ][3]<= -18; ws[4][4 ][4]<=-200; ws[4][4 ][5]<=-269; ws[4][4 ][6]<=-138; ws[4][4 ][7]<=  32; ws[4][4 ][8]<= 115; ws[4][4 ][9]<= 140; ws[4][4 ][10]<= 106; ws[4][4 ][11]<=-177; ws[4][4 ][12]<=-271; ws[4][4 ][13]<=-162; ws[4][4 ][14]<=  15; ws[4][4 ][15]<=  23; ws[4][4 ][16]<= 123; ws[4][4 ][17]<=  87; ws[4][4 ][18]<= -72; ws[4][4 ][19]<=-184; ws[4][4 ][20]<=-157; ws[4][4 ][21]<=  32; ws[4][4 ][22]<= -45; ws[4][4 ][23]<=   8; ws[4][4 ][24]<= 123; ws[4][4 ][25]<=  56; ws[4][4 ][26]<= -24; ws[4][4 ][27]<= -28; ws[4][4 ][28]<=  42; ws[4][4 ][29]<= -60; ws[4][4 ][30]<=-134; ws[4][4 ][31]<=  40; ws[4][4 ][32]<= 142; ws[4][4 ][33]<= 154; ws[4][4 ][34]<=  45; ws[4][4 ][35]<=  48; ws[4][4 ][36]<= -57; ws[4][4 ][37]<=-127; ws[4][4 ][38]<= -45; ws[4][4 ][39]<= 187; ws[4][4 ][40]<= 199; ws[4][4 ][41]<= 142; ws[4][4 ][42]<=  37; ws[4][4 ][43]<= -12; ws[4][4 ][44]<= -93; ws[4][4 ][45]<=-123; ws[4][4 ][46]<=  87; ws[4][4 ][47]<= 268; ws[4][4 ][48]<= 245;
        ws[4][5 ][0]<=  64; ws[4][5 ][1]<= 112; ws[4][5 ][2]<= 109; ws[4][5 ][3]<= -25; ws[4][5 ][4]<=-115; ws[4][5 ][5]<=-104; ws[4][5 ][6]<=  85; ws[4][5 ][7]<=  92; ws[4][5 ][8]<= 139; ws[4][5 ][9]<=  55; ws[4][5 ][10]<=  14; ws[4][5 ][11]<= -81; ws[4][5 ][12]<= -45; ws[4][5 ][13]<=  58; ws[4][5 ][14]<=  85; ws[4][5 ][15]<= 104; ws[4][5 ][16]<=  57; ws[4][5 ][17]<= 123; ws[4][5 ][18]<=  37; ws[4][5 ][19]<= -19; ws[4][5 ][20]<=  80; ws[4][5 ][21]<=  29; ws[4][5 ][22]<=  59; ws[4][5 ][23]<=  90; ws[4][5 ][24]<= 125; ws[4][5 ][25]<= 115; ws[4][5 ][26]<=  32; ws[4][5 ][27]<= 112; ws[4][5 ][28]<= -20; ws[4][5 ][29]<=   2; ws[4][5 ][30]<=  45; ws[4][5 ][31]<= 121; ws[4][5 ][32]<= 112; ws[4][5 ][33]<= 112; ws[4][5 ][34]<= 127; ws[4][5 ][35]<= -21; ws[4][5 ][36]<= -66; ws[4][5 ][37]<= -52; ws[4][5 ][38]<=  97; ws[4][5 ][39]<= 142; ws[4][5 ][40]<= 160; ws[4][5 ][41]<= 178; ws[4][5 ][42]<=-109; ws[4][5 ][43]<= -71; ws[4][5 ][44]<=   0; ws[4][5 ][45]<=  60; ws[4][5 ][46]<= 105; ws[4][5 ][47]<= 189; ws[4][5 ][48]<= 185;
        ws[4][6 ][0]<= 136; ws[4][6 ][1]<=  11; ws[4][6 ][2]<= -64; ws[4][6 ][3]<=  57; ws[4][6 ][4]<=  40; ws[4][6 ][5]<=-113; ws[4][6 ][6]<=-224; ws[4][6 ][7]<=  81; ws[4][6 ][8]<=  21; ws[4][6 ][9]<= -20; ws[4][6 ][10]<=  55; ws[4][6 ][11]<=  34; ws[4][6 ][12]<=-126; ws[4][6 ][13]<=-209; ws[4][6 ][14]<=  99; ws[4][6 ][15]<=  72; ws[4][6 ][16]<= -57; ws[4][6 ][17]<=  87; ws[4][6 ][18]<=  20; ws[4][6 ][19]<= -59; ws[4][6 ][20]<=-174; ws[4][6 ][21]<=  59; ws[4][6 ][22]<=  18; ws[4][6 ][23]<=   1; ws[4][6 ][24]<= 101; ws[4][6 ][25]<= 103; ws[4][6 ][26]<= -42; ws[4][6 ][27]<=-127; ws[4][6 ][28]<=  33; ws[4][6 ][29]<=   6; ws[4][6 ][30]<= -81; ws[4][6 ][31]<= 101; ws[4][6 ][32]<= 117; ws[4][6 ][33]<= -30; ws[4][6 ][34]<=-159; ws[4][6 ][35]<=  99; ws[4][6 ][36]<=-105; ws[4][6 ][37]<=-100; ws[4][6 ][38]<=  34; ws[4][6 ][39]<=  65; ws[4][6 ][40]<=  12; ws[4][6 ][41]<=-103; ws[4][6 ][42]<=  71; ws[4][6 ][43]<= -97; ws[4][6 ][44]<=-186; ws[4][6 ][45]<= -46; ws[4][6 ][46]<=  20; ws[4][6 ][47]<= -19; ws[4][6 ][48]<=-110;
        ws[4][7 ][0]<= -24; ws[4][7 ][1]<=  13; ws[4][7 ][2]<=  18; ws[4][7 ][3]<=  18; ws[4][7 ][4]<=  85; ws[4][7 ][5]<=  64; ws[4][7 ][6]<=  49; ws[4][7 ][7]<= -44; ws[4][7 ][8]<= -33; ws[4][7 ][9]<=   6; ws[4][7 ][10]<=  79; ws[4][7 ][11]<=  64; ws[4][7 ][12]<=  88; ws[4][7 ][13]<=  45; ws[4][7 ][14]<= -86; ws[4][7 ][15]<=  -8; ws[4][7 ][16]<=  -1; ws[4][7 ][17]<= 115; ws[4][7 ][18]<=  90; ws[4][7 ][19]<= 152; ws[4][7 ][20]<=  64; ws[4][7 ][21]<= -15; ws[4][7 ][22]<=  25; ws[4][7 ][23]<=  61; ws[4][7 ][24]<=  71; ws[4][7 ][25]<= 143; ws[4][7 ][26]<= 159; ws[4][7 ][27]<= 116; ws[4][7 ][28]<=  60; ws[4][7 ][29]<= 114; ws[4][7 ][30]<=  53; ws[4][7 ][31]<=  84; ws[4][7 ][32]<=  67; ws[4][7 ][33]<= 128; ws[4][7 ][34]<= 155; ws[4][7 ][35]<=  58; ws[4][7 ][36]<= 115; ws[4][7 ][37]<=  77; ws[4][7 ][38]<=  70; ws[4][7 ][39]<= 120; ws[4][7 ][40]<= 128; ws[4][7 ][41]<= 184; ws[4][7 ][42]<=  46; ws[4][7 ][43]<= 114; ws[4][7 ][44]<=  34; ws[4][7 ][45]<=  15; ws[4][7 ][46]<=  57; ws[4][7 ][47]<= 196; ws[4][7 ][48]<= 205;
        ws[4][8 ][0]<=  18; ws[4][8 ][1]<= -93; ws[4][8 ][2]<= -27; ws[4][8 ][3]<=   1; ws[4][8 ][4]<= -33; ws[4][8 ][5]<=-107; ws[4][8 ][6]<= -46; ws[4][8 ][7]<=  71; ws[4][8 ][8]<= -42; ws[4][8 ][9]<=  12; ws[4][8 ][10]<=   0; ws[4][8 ][11]<= -17; ws[4][8 ][12]<= -88; ws[4][8 ][13]<= -98; ws[4][8 ][14]<= 103; ws[4][8 ][15]<=  32; ws[4][8 ][16]<=  18; ws[4][8 ][17]<=  81; ws[4][8 ][18]<=  75; ws[4][8 ][19]<= -31; ws[4][8 ][20]<= -89; ws[4][8 ][21]<=  89; ws[4][8 ][22]<= -16; ws[4][8 ][23]<=  27; ws[4][8 ][24]<=  26; ws[4][8 ][25]<= 131; ws[4][8 ][26]<=  21; ws[4][8 ][27]<=  20; ws[4][8 ][28]<=  26; ws[4][8 ][29]<= -16; ws[4][8 ][30]<= -33; ws[4][8 ][31]<=  31; ws[4][8 ][32]<= 139; ws[4][8 ][33]<=  56; ws[4][8 ][34]<=  56; ws[4][8 ][35]<=   4; ws[4][8 ][36]<= -41; ws[4][8 ][37]<=-101; ws[4][8 ][38]<=  52; ws[4][8 ][39]<= 208; ws[4][8 ][40]<= 213; ws[4][8 ][41]<= 162; ws[4][8 ][42]<= -66; ws[4][8 ][43]<= -78; ws[4][8 ][44]<= -52; ws[4][8 ][45]<=  12; ws[4][8 ][46]<= 188; ws[4][8 ][47]<= 194; ws[4][8 ][48]<= 207;
        ws[4][9 ][0]<=  91; ws[4][9 ][1]<= 108; ws[4][9 ][2]<= -65; ws[4][9 ][3]<= -91; ws[4][9 ][4]<= -35; ws[4][9 ][5]<=  55; ws[4][9 ][6]<=  26; ws[4][9 ][7]<=  59; ws[4][9 ][8]<=  56; ws[4][9 ][9]<= -32; ws[4][9 ][10]<=-104; ws[4][9 ][11]<= -56; ws[4][9 ][12]<=  13; ws[4][9 ][13]<= -34; ws[4][9 ][14]<=   3; ws[4][9 ][15]<=   3; ws[4][9 ][16]<= -34; ws[4][9 ][17]<= -60; ws[4][9 ][18]<= -75; ws[4][9 ][19]<=  45; ws[4][9 ][20]<= -45; ws[4][9 ][21]<=  48; ws[4][9 ][22]<=  -4; ws[4][9 ][23]<= -34; ws[4][9 ][24]<=-135; ws[4][9 ][25]<= -89; ws[4][9 ][26]<=  -3; ws[4][9 ][27]<= -11; ws[4][9 ][28]<=  56; ws[4][9 ][29]<=  41; ws[4][9 ][30]<=  20; ws[4][9 ][31]<=-119; ws[4][9 ][32]<=-125; ws[4][9 ][33]<= -74; ws[4][9 ][34]<= -38; ws[4][9 ][35]<=  91; ws[4][9 ][36]<=  60; ws[4][9 ][37]<=   5; ws[4][9 ][38]<=-128; ws[4][9 ][39]<=-142; ws[4][9 ][40]<= -94; ws[4][9 ][41]<=  59; ws[4][9 ][42]<= 153; ws[4][9 ][43]<=  87; ws[4][9 ][44]<=  34; ws[4][9 ][45]<= -79; ws[4][9 ][46]<=-188; ws[4][9 ][47]<=-102; ws[4][9 ][48]<=   7;
        ws[4][10][0]<= 118; ws[4][10][1]<=  39; ws[4][10][2]<= -47; ws[4][10][3]<= -77; ws[4][10][4]<=  35; ws[4][10][5]<=  83; ws[4][10][6]<= 188; ws[4][10][7]<=  77; ws[4][10][8]<=  65; ws[4][10][9]<=  26; ws[4][10][10]<= -54; ws[4][10][11]<=   8; ws[4][10][12]<= 112; ws[4][10][13]<= 211; ws[4][10][14]<=  58; ws[4][10][15]<=  48; ws[4][10][16]<=  34; ws[4][10][17]<=  40; ws[4][10][18]<=  10; ws[4][10][19]<=  86; ws[4][10][20]<= 187; ws[4][10][21]<=  -5; ws[4][10][22]<=  65; ws[4][10][23]<=  39; ws[4][10][24]<=   6; ws[4][10][25]<=  40; ws[4][10][26]<=  70; ws[4][10][27]<= 180; ws[4][10][28]<=  31; ws[4][10][29]<=  13; ws[4][10][30]<= -13; ws[4][10][31]<=  39; ws[4][10][32]<=  83; ws[4][10][33]<= 104; ws[4][10][34]<=  54; ws[4][10][35]<= -34; ws[4][10][36]<= -17; ws[4][10][37]<= -67; ws[4][10][38]<= -80; ws[4][10][39]<=  64; ws[4][10][40]<=  70; ws[4][10][41]<=  58; ws[4][10][42]<= -36; ws[4][10][43]<= -63; ws[4][10][44]<=-197; ws[4][10][45]<=-120; ws[4][10][46]<=  -7; ws[4][10][47]<= 100; ws[4][10][48]<= 115;
        ws[4][11][0]<=-107; ws[4][11][1]<= 137; ws[4][11][2]<= 197; ws[4][11][3]<= 108; ws[4][11][4]<=  79; ws[4][11][5]<=  30; ws[4][11][6]<= -32; ws[4][11][7]<= -77; ws[4][11][8]<= 112; ws[4][11][9]<= 137; ws[4][11][10]<= 139; ws[4][11][11]<=  64; ws[4][11][12]<= -22; ws[4][11][13]<= -83; ws[4][11][14]<=-126; ws[4][11][15]<=  20; ws[4][11][16]<= 128; ws[4][11][17]<=  85; ws[4][11][18]<= -10; ws[4][11][19]<= -80; ws[4][11][20]<= -41; ws[4][11][21]<= -81; ws[4][11][22]<= -19; ws[4][11][23]<= 130; ws[4][11][24]<=  83; ws[4][11][25]<=  24; ws[4][11][26]<= -67; ws[4][11][27]<= -85; ws[4][11][28]<= -94; ws[4][11][29]<=  23; ws[4][11][30]<=  92; ws[4][11][31]<=  81; ws[4][11][32]<=  -6; ws[4][11][33]<= -93; ws[4][11][34]<= -23; ws[4][11][35]<= -98; ws[4][11][36]<= -55; ws[4][11][37]<=  71; ws[4][11][38]<=  64; ws[4][11][39]<=   9; ws[4][11][40]<= -34; ws[4][11][41]<= 152; ws[4][11][42]<= -87; ws[4][11][43]<=-115; ws[4][11][44]<=  63; ws[4][11][45]<=  56; ws[4][11][46]<=  20; ws[4][11][47]<=  17; ws[4][11][48]<= 289;
        ws[4][12][0]<= 125; ws[4][12][1]<=  99; ws[4][12][2]<= 128; ws[4][12][3]<= 122; ws[4][12][4]<=  88; ws[4][12][5]<= 159; ws[4][12][6]<= 141; ws[4][12][7]<=  77; ws[4][12][8]<= 109; ws[4][12][9]<=  83; ws[4][12][10]<=  33; ws[4][12][11]<=  26; ws[4][12][12]<=  80; ws[4][12][13]<= 129; ws[4][12][14]<=  43; ws[4][12][15]<=  45; ws[4][12][16]<=  31; ws[4][12][17]<=   2; ws[4][12][18]<= -50; ws[4][12][19]<= -29; ws[4][12][20]<= 128; ws[4][12][21]<=  15; ws[4][12][22]<=  87; ws[4][12][23]<=  33; ws[4][12][24]<=  59; ws[4][12][25]<= -27; ws[4][12][26]<=  -5; ws[4][12][27]<= 103; ws[4][12][28]<=   2; ws[4][12][29]<=  -2; ws[4][12][30]<=  50; ws[4][12][31]<=  -4; ws[4][12][32]<= -30; ws[4][12][33]<= -17; ws[4][12][34]<=  57; ws[4][12][35]<=-137; ws[4][12][36]<= -50; ws[4][12][37]<=   0; ws[4][12][38]<= -10; ws[4][12][39]<= -28; ws[4][12][40]<= -14; ws[4][12][41]<=  85; ws[4][12][42]<=-162; ws[4][12][43]<=-112; ws[4][12][44]<= -81; ws[4][12][45]<=  40; ws[4][12][46]<= -38; ws[4][12][47]<=   0; ws[4][12][48]<=  40;
        ws[4][13][0]<= -43; ws[4][13][1]<=  11; ws[4][13][2]<= 138; ws[4][13][3]<= 131; ws[4][13][4]<=  62; ws[4][13][5]<= -11; ws[4][13][6]<= -30; ws[4][13][7]<=  18; ws[4][13][8]<=  29; ws[4][13][9]<= 127; ws[4][13][10]<= 136; ws[4][13][11]<= 114; ws[4][13][12]<=  -4; ws[4][13][13]<= -58; ws[4][13][14]<= -21; ws[4][13][15]<=  16; ws[4][13][16]<= 139; ws[4][13][17]<= 175; ws[4][13][18]<= 119; ws[4][13][19]<= -17; ws[4][13][20]<=-100; ws[4][13][21]<=   7; ws[4][13][22]<=  13; ws[4][13][23]<=  91; ws[4][13][24]<= 171; ws[4][13][25]<= 109; ws[4][13][26]<= -86; ws[4][13][27]<=-125; ws[4][13][28]<= -19; ws[4][13][29]<= -14; ws[4][13][30]<= 101; ws[4][13][31]<= 197; ws[4][13][32]<= 104; ws[4][13][33]<= -74; ws[4][13][34]<= -60; ws[4][13][35]<= -86; ws[4][13][36]<=-117; ws[4][13][37]<=  79; ws[4][13][38]<= 132; ws[4][13][39]<=  50; ws[4][13][40]<= -93; ws[4][13][41]<= -53; ws[4][13][42]<=-202; ws[4][13][43]<= -87; ws[4][13][44]<=   9; ws[4][13][45]<= 102; ws[4][13][46]<=  22; ws[4][13][47]<= -99; ws[4][13][48]<= -54;
        ws[4][14][0]<=  -1; ws[4][14][1]<= -78; ws[4][14][2]<= -29; ws[4][14][3]<= -51; ws[4][14][4]<= -64; ws[4][14][5]<= -97; ws[4][14][6]<=-144; ws[4][14][7]<= -62; ws[4][14][8]<=-105; ws[4][14][9]<=  -4; ws[4][14][10]<=  22; ws[4][14][11]<= -39; ws[4][14][12]<= -55; ws[4][14][13]<= -87; ws[4][14][14]<= -26; ws[4][14][15]<= -96; ws[4][14][16]<= -53; ws[4][14][17]<=  86; ws[4][14][18]<=  87; ws[4][14][19]<=   9; ws[4][14][20]<=  -7; ws[4][14][21]<=  35; ws[4][14][22]<= -76; ws[4][14][23]<=  26; ws[4][14][24]<=  55; ws[4][14][25]<=  53; ws[4][14][26]<= 101; ws[4][14][27]<=  53; ws[4][14][28]<=  18; ws[4][14][29]<= -54; ws[4][14][30]<= -38; ws[4][14][31]<= 106; ws[4][14][32]<=  82; ws[4][14][33]<= 121; ws[4][14][34]<= 140; ws[4][14][35]<= 109; ws[4][14][36]<=  -6; ws[4][14][37]<= -27; ws[4][14][38]<=  58; ws[4][14][39]<= 108; ws[4][14][40]<= 158; ws[4][14][41]<= 123; ws[4][14][42]<=  89; ws[4][14][43]<=  49; ws[4][14][44]<=  32; ws[4][14][45]<=  22; ws[4][14][46]<= 109; ws[4][14][47]<=  92; ws[4][14][48]<= 191;
        ws[4][15][0]<= 134; ws[4][15][1]<= 133; ws[4][15][2]<= 106; ws[4][15][3]<=  85; ws[4][15][4]<= 138; ws[4][15][5]<= 121; ws[4][15][6]<=  18; ws[4][15][7]<=  24; ws[4][15][8]<=  85; ws[4][15][9]<= 107; ws[4][15][10]<=  48; ws[4][15][11]<= 132; ws[4][15][12]<= 148; ws[4][15][13]<=  11; ws[4][15][14]<=   8; ws[4][15][15]<=  16; ws[4][15][16]<=  93; ws[4][15][17]<=  21; ws[4][15][18]<=  23; ws[4][15][19]<= 106; ws[4][15][20]<=  -8; ws[4][15][21]<= -40; ws[4][15][22]<=  74; ws[4][15][23]<=  90; ws[4][15][24]<=  60; ws[4][15][25]<= -50; ws[4][15][26]<=   5; ws[4][15][27]<=  17; ws[4][15][28]<= -31; ws[4][15][29]<=  45; ws[4][15][30]<= 102; ws[4][15][31]<= -37; ws[4][15][32]<=-133; ws[4][15][33]<= -84; ws[4][15][34]<= -28; ws[4][15][35]<=  36; ws[4][15][36]<=  45; ws[4][15][37]<= 110; ws[4][15][38]<= -17; ws[4][15][39]<=-145; ws[4][15][40]<=-180; ws[4][15][41]<=-147; ws[4][15][42]<=  51; ws[4][15][43]<=  -1; ws[4][15][44]<=  10; ws[4][15][45]<=-132; ws[4][15][46]<=-250; ws[4][15][47]<=-198; ws[4][15][48]<=-176;

        ws[5][0 ][0]<=  48; ws[5][0 ][1]<= -47; ws[5][0 ][2]<= -34; ws[5][0 ][3]<=  52; ws[5][0 ][4]<= 145; ws[5][0 ][5]<=  24; ws[5][0 ][6]<= -55; ws[5][0 ][7]<= 196; ws[5][0 ][8]<= 107; ws[5][0 ][9]<=  56; ws[5][0 ][10]<=  87; ws[5][0 ][11]<=  51; ws[5][0 ][12]<= -12; ws[5][0 ][13]<=-108; ws[5][0 ][14]<= 212; ws[5][0 ][15]<= 162; ws[5][0 ][16]<=  34; ws[5][0 ][17]<= -80; ws[5][0 ][18]<= -42; ws[5][0 ][19]<= -21; ws[5][0 ][20]<= -46; ws[5][0 ][21]<= 146; ws[5][0 ][22]<=  57; ws[5][0 ][23]<= -50; ws[5][0 ][24]<=-156; ws[5][0 ][25]<= -17; ws[5][0 ][26]<=  37; ws[5][0 ][27]<= -36; ws[5][0 ][28]<=   1; ws[5][0 ][29]<=  28; ws[5][0 ][30]<= -84; ws[5][0 ][31]<=-189; ws[5][0 ][32]<= -75; ws[5][0 ][33]<= 108; ws[5][0 ][34]<= -48; ws[5][0 ][35]<=-116; ws[5][0 ][36]<= -85; ws[5][0 ][37]<=   2; ws[5][0 ][38]<=-150; ws[5][0 ][39]<= -97; ws[5][0 ][40]<=  65; ws[5][0 ][41]<=-113; ws[5][0 ][42]<=-142; ws[5][0 ][43]<=  41; ws[5][0 ][44]<= 152; ws[5][0 ][45]<= -38; ws[5][0 ][46]<=-128; ws[5][0 ][47]<= -12; ws[5][0 ][48]<=-102;
        ws[5][1 ][0]<= 156; ws[5][1 ][1]<= -63; ws[5][1 ][2]<=-145; ws[5][1 ][3]<=-176; ws[5][1 ][4]<=-221; ws[5][1 ][5]<=-194; ws[5][1 ][6]<=-285; ws[5][1 ][7]<= -58; ws[5][1 ][8]<=-168; ws[5][1 ][9]<=-162; ws[5][1 ][10]<=-104; ws[5][1 ][11]<= -72; ws[5][1 ][12]<= -64; ws[5][1 ][13]<=-237; ws[5][1 ][14]<=-155; ws[5][1 ][15]<= -74; ws[5][1 ][16]<= -58; ws[5][1 ][17]<=   0; ws[5][1 ][18]<= -31; ws[5][1 ][19]<=  -2; ws[5][1 ][20]<=-161; ws[5][1 ][21]<= -66; ws[5][1 ][22]<=   1; ws[5][1 ][23]<= -70; ws[5][1 ][24]<=  -4; ws[5][1 ][25]<=  12; ws[5][1 ][26]<= -21; ws[5][1 ][27]<=-185; ws[5][1 ][28]<= -39; ws[5][1 ][29]<= -29; ws[5][1 ][30]<=  37; ws[5][1 ][31]<=   7; ws[5][1 ][32]<= -28; ws[5][1 ][33]<= -91; ws[5][1 ][34]<=-150; ws[5][1 ][35]<= -92; ws[5][1 ][36]<= -71; ws[5][1 ][37]<= -41; ws[5][1 ][38]<=  -6; ws[5][1 ][39]<= -91; ws[5][1 ][40]<= -43; ws[5][1 ][41]<=-188; ws[5][1 ][42]<=-229; ws[5][1 ][43]<=-228; ws[5][1 ][44]<=-108; ws[5][1 ][45]<= -92; ws[5][1 ][46]<=-116; ws[5][1 ][47]<=-144; ws[5][1 ][48]<=-287;
        ws[5][2 ][0]<= -88; ws[5][2 ][1]<=-136; ws[5][2 ][2]<=-157; ws[5][2 ][3]<=-173; ws[5][2 ][4]<=-111; ws[5][2 ][5]<= -70; ws[5][2 ][6]<=-135; ws[5][2 ][7]<= -44; ws[5][2 ][8]<= -37; ws[5][2 ][9]<=-105; ws[5][2 ][10]<= -76; ws[5][2 ][11]<=-133; ws[5][2 ][12]<= -34; ws[5][2 ][13]<= -81; ws[5][2 ][14]<= -16; ws[5][2 ][15]<=-113; ws[5][2 ][16]<= -25; ws[5][2 ][17]<= -94; ws[5][2 ][18]<= -67; ws[5][2 ][19]<= -69; ws[5][2 ][20]<= -29; ws[5][2 ][21]<= -95; ws[5][2 ][22]<=-113; ws[5][2 ][23]<= -98; ws[5][2 ][24]<=   1; ws[5][2 ][25]<= -51; ws[5][2 ][26]<=  17; ws[5][2 ][27]<= -31; ws[5][2 ][28]<= -30; ws[5][2 ][29]<=-129; ws[5][2 ][30]<= -34; ws[5][2 ][31]<= -13; ws[5][2 ][32]<= -19; ws[5][2 ][33]<=  15; ws[5][2 ][34]<=  73; ws[5][2 ][35]<=  -9; ws[5][2 ][36]<= -55; ws[5][2 ][37]<= -91; ws[5][2 ][38]<=  60; ws[5][2 ][39]<=   4; ws[5][2 ][40]<=  60; ws[5][2 ][41]<=  68; ws[5][2 ][42]<=  -5; ws[5][2 ][43]<= -25; ws[5][2 ][44]<= -96; ws[5][2 ][45]<=  32; ws[5][2 ][46]<= 132; ws[5][2 ][47]<= 125; ws[5][2 ][48]<= 120;
        ws[5][3 ][0]<= -89; ws[5][3 ][1]<= -17; ws[5][3 ][2]<=  78; ws[5][3 ][3]<=  88; ws[5][3 ][4]<=  41; ws[5][3 ][5]<=  28; ws[5][3 ][6]<=  82; ws[5][3 ][7]<= -74; ws[5][3 ][8]<=  50; ws[5][3 ][9]<= 119; ws[5][3 ][10]<= 125; ws[5][3 ][11]<= -11; ws[5][3 ][12]<= -37; ws[5][3 ][13]<=  25; ws[5][3 ][14]<= -85; ws[5][3 ][15]<=  39; ws[5][3 ][16]<=  98; ws[5][3 ][17]<= 170; ws[5][3 ][18]<=  60; ws[5][3 ][19]<=   5; ws[5][3 ][20]<=  -9; ws[5][3 ][21]<= -81; ws[5][3 ][22]<= -39; ws[5][3 ][23]<= 138; ws[5][3 ][24]<= 134; ws[5][3 ][25]<=  44; ws[5][3 ][26]<=  15; ws[5][3 ][27]<=  30; ws[5][3 ][28]<=  47; ws[5][3 ][29]<=  -2; ws[5][3 ][30]<=  20; ws[5][3 ][31]<=  88; ws[5][3 ][32]<=  84; ws[5][3 ][33]<=   8; ws[5][3 ][34]<=  29; ws[5][3 ][35]<=  80; ws[5][3 ][36]<=  31; ws[5][3 ][37]<=  20; ws[5][3 ][38]<= 139; ws[5][3 ][39]<= 116; ws[5][3 ][40]<=  30; ws[5][3 ][41]<=  45; ws[5][3 ][42]<= 105; ws[5][3 ][43]<=  19; ws[5][3 ][44]<=  39; ws[5][3 ][45]<= 155; ws[5][3 ][46]<=  97; ws[5][3 ][47]<=  64; ws[5][3 ][48]<=   8;
        ws[5][4 ][0]<=-101; ws[5][4 ][1]<= -34; ws[5][4 ][2]<=   1; ws[5][4 ][3]<=  60; ws[5][4 ][4]<=  67; ws[5][4 ][5]<=  68; ws[5][4 ][6]<=  45; ws[5][4 ][7]<= -71; ws[5][4 ][8]<= -50; ws[5][4 ][9]<= -58; ws[5][4 ][10]<=  44; ws[5][4 ][11]<=  50; ws[5][4 ][12]<=  70; ws[5][4 ][13]<=  34; ws[5][4 ][14]<=  27; ws[5][4 ][15]<= -27; ws[5][4 ][16]<= -83; ws[5][4 ][17]<= -13; ws[5][4 ][18]<=  40; ws[5][4 ][19]<=  25; ws[5][4 ][20]<=  90; ws[5][4 ][21]<=  16; ws[5][4 ][22]<=   2; ws[5][4 ][23]<=  -9; ws[5][4 ][24]<=  39; ws[5][4 ][25]<=  65; ws[5][4 ][26]<=  60; ws[5][4 ][27]<=  54; ws[5][4 ][28]<=  85; ws[5][4 ][29]<=  28; ws[5][4 ][30]<= -14; ws[5][4 ][31]<=  64; ws[5][4 ][32]<= 110; ws[5][4 ][33]<= 114; ws[5][4 ][34]<= 122; ws[5][4 ][35]<= 140; ws[5][4 ][36]<=  31; ws[5][4 ][37]<= -27; ws[5][4 ][38]<=  38; ws[5][4 ][39]<=  66; ws[5][4 ][40]<=  94; ws[5][4 ][41]<= 107; ws[5][4 ][42]<= 156; ws[5][4 ][43]<=  76; ws[5][4 ][44]<= -39; ws[5][4 ][45]<=   3; ws[5][4 ][46]<= 130; ws[5][4 ][47]<=  96; ws[5][4 ][48]<= 180;
        ws[5][5 ][0]<= 148; ws[5][5 ][1]<=  87; ws[5][5 ][2]<= 109; ws[5][5 ][3]<= 164; ws[5][5 ][4]<=  62; ws[5][5 ][5]<= -17; ws[5][5 ][6]<=  77; ws[5][5 ][7]<= 105; ws[5][5 ][8]<=  69; ws[5][5 ][9]<=  38; ws[5][5 ][10]<= 128; ws[5][5 ][11]<=  70; ws[5][5 ][12]<=   9; ws[5][5 ][13]<= -39; ws[5][5 ][14]<=  13; ws[5][5 ][15]<= -15; ws[5][5 ][16]<=  17; ws[5][5 ][17]<=  68; ws[5][5 ][18]<=  61; ws[5][5 ][19]<= -30; ws[5][5 ][20]<=  -7; ws[5][5 ][21]<=  31; ws[5][5 ][22]<=  45; ws[5][5 ][23]<= -15; ws[5][5 ][24]<= 100; ws[5][5 ][25]<=  50; ws[5][5 ][26]<= -55; ws[5][5 ][27]<= -50; ws[5][5 ][28]<=  28; ws[5][5 ][29]<=  18; ws[5][5 ][30]<=  73; ws[5][5 ][31]<=   9; ws[5][5 ][32]<= -28; ws[5][5 ][33]<= -90; ws[5][5 ][34]<= -92; ws[5][5 ][35]<=  27; ws[5][5 ][36]<=  98; ws[5][5 ][37]<=  24; ws[5][5 ][38]<=  11; ws[5][5 ][39]<= -62; ws[5][5 ][40]<=-110; ws[5][5 ][41]<=-123; ws[5][5 ][42]<= 135; ws[5][5 ][43]<= 172; ws[5][5 ][44]<= 120; ws[5][5 ][45]<=  27; ws[5][5 ][46]<=-107; ws[5][5 ][47]<= -76; ws[5][5 ][48]<=-107;
        ws[5][6 ][0]<= -71; ws[5][6 ][1]<= -31; ws[5][6 ][2]<= -91; ws[5][6 ][3]<= -24; ws[5][6 ][4]<=  31; ws[5][6 ][5]<= 172; ws[5][6 ][6]<=-111; ws[5][6 ][7]<= -23; ws[5][6 ][8]<= -64; ws[5][6 ][9]<=   5; ws[5][6 ][10]<= -11; ws[5][6 ][11]<= 104; ws[5][6 ][12]<= 219; ws[5][6 ][13]<= -94; ws[5][6 ][14]<= -65; ws[5][6 ][15]<=-114; ws[5][6 ][16]<= -57; ws[5][6 ][17]<= -54; ws[5][6 ][18]<= 156; ws[5][6 ][19]<= 278; ws[5][6 ][20]<= -35; ws[5][6 ][21]<= -70; ws[5][6 ][22]<=-153; ws[5][6 ][23]<= -92; ws[5][6 ][24]<= -11; ws[5][6 ][25]<= 157; ws[5][6 ][26]<= 242; ws[5][6 ][27]<= -31; ws[5][6 ][28]<= -51; ws[5][6 ][29]<=-130; ws[5][6 ][30]<= -49; ws[5][6 ][31]<=  46; ws[5][6 ][32]<= 147; ws[5][6 ][33]<= 127; ws[5][6 ][34]<=-175; ws[5][6 ][35]<= 106; ws[5][6 ][36]<=  -2; ws[5][6 ][37]<=  35; ws[5][6 ][38]<=  52; ws[5][6 ][39]<= 123; ws[5][6 ][40]<=  -8; ws[5][6 ][41]<=-168; ws[5][6 ][42]<= 186; ws[5][6 ][43]<=  57; ws[5][6 ][44]<=  84; ws[5][6 ][45]<=  85; ws[5][6 ][46]<=  43; ws[5][6 ][47]<= -34; ws[5][6 ][48]<=   2;
        ws[5][7 ][0]<=-110; ws[5][7 ][1]<=  66; ws[5][7 ][2]<= 107; ws[5][7 ][3]<=-140; ws[5][7 ][4]<=-120; ws[5][7 ][5]<= -79; ws[5][7 ][6]<= -89; ws[5][7 ][7]<= -64; ws[5][7 ][8]<=  83; ws[5][7 ][9]<=  95; ws[5][7 ][10]<= -93; ws[5][7 ][11]<= -64; ws[5][7 ][12]<=  -8; ws[5][7 ][13]<= -39; ws[5][7 ][14]<= -64; ws[5][7 ][15]<= 102; ws[5][7 ][16]<= 118; ws[5][7 ][17]<= -47; ws[5][7 ][18]<= -75; ws[5][7 ][19]<=  60; ws[5][7 ][20]<=  31; ws[5][7 ][21]<=-152; ws[5][7 ][22]<=  65; ws[5][7 ][23]<= 129; ws[5][7 ][24]<= -40; ws[5][7 ][25]<= -50; ws[5][7 ][26]<= 110; ws[5][7 ][27]<=  72; ws[5][7 ][28]<=-106; ws[5][7 ][29]<=  24; ws[5][7 ][30]<= 145; ws[5][7 ][31]<= -67; ws[5][7 ][32]<= -59; ws[5][7 ][33]<= 153; ws[5][7 ][34]<=  79; ws[5][7 ][35]<= -31; ws[5][7 ][36]<= 105; ws[5][7 ][37]<= 192; ws[5][7 ][38]<= -64; ws[5][7 ][39]<= -19; ws[5][7 ][40]<=  58; ws[5][7 ][41]<= 164; ws[5][7 ][42]<=  64; ws[5][7 ][43]<= 143; ws[5][7 ][44]<= 251; ws[5][7 ][45]<=  51; ws[5][7 ][46]<= -32; ws[5][7 ][47]<= 103; ws[5][7 ][48]<= 132;
        ws[5][8 ][0]<= -24; ws[5][8 ][1]<= 237; ws[5][8 ][2]<= 129; ws[5][8 ][3]<= -64; ws[5][8 ][4]<= -85; ws[5][8 ][5]<= -31; ws[5][8 ][6]<= 120; ws[5][8 ][7]<= -43; ws[5][8 ][8]<= 157; ws[5][8 ][9]<= 148; ws[5][8 ][10]<=  13; ws[5][8 ][11]<= -44; ws[5][8 ][12]<= -31; ws[5][8 ][13]<= 119; ws[5][8 ][14]<=-136; ws[5][8 ][15]<= 149; ws[5][8 ][16]<= 105; ws[5][8 ][17]<=   7; ws[5][8 ][18]<= -22; ws[5][8 ][19]<=  15; ws[5][8 ][20]<= 121; ws[5][8 ][21]<=-156; ws[5][8 ][22]<=  38; ws[5][8 ][23]<= 133; ws[5][8 ][24]<= -39; ws[5][8 ][25]<=  10; ws[5][8 ][26]<= -14; ws[5][8 ][27]<= 192; ws[5][8 ][28]<=-146; ws[5][8 ][29]<=  17; ws[5][8 ][30]<=  27; ws[5][8 ][31]<=  15; ws[5][8 ][32]<= -80; ws[5][8 ][33]<=  -2; ws[5][8 ][34]<= 167; ws[5][8 ][35]<=-131; ws[5][8 ][36]<= -58; ws[5][8 ][37]<=  -2; ws[5][8 ][38]<= -69; ws[5][8 ][39]<= -55; ws[5][8 ][40]<=   0; ws[5][8 ][41]<= 183; ws[5][8 ][42]<= -31; ws[5][8 ][43]<= -68; ws[5][8 ][44]<= -85; ws[5][8 ][45]<=-117; ws[5][8 ][46]<=-100; ws[5][8 ][47]<=  16; ws[5][8 ][48]<= 178;
        ws[5][9 ][0]<= -66; ws[5][9 ][1]<= -67; ws[5][9 ][2]<=  75; ws[5][9 ][3]<= 133; ws[5][9 ][4]<= 122; ws[5][9 ][5]<=  46; ws[5][9 ][6]<=-168; ws[5][9 ][7]<=-167; ws[5][9 ][8]<=-154; ws[5][9 ][9]<=  70; ws[5][9 ][10]<= 115; ws[5][9 ][11]<= 175; ws[5][9 ][12]<= 143; ws[5][9 ][13]<= -96; ws[5][9 ][14]<= -55; ws[5][9 ][15]<= -63; ws[5][9 ][16]<= 100; ws[5][9 ][17]<= 106; ws[5][9 ][18]<=  75; ws[5][9 ][19]<= 118; ws[5][9 ][20]<= -83; ws[5][9 ][21]<=  41; ws[5][9 ][22]<=  30; ws[5][9 ][23]<= 115; ws[5][9 ][24]<=  -2; ws[5][9 ][25]<=  38; ws[5][9 ][26]<= 107; ws[5][9 ][27]<= -53; ws[5][9 ][28]<=  26; ws[5][9 ][29]<=  -5; ws[5][9 ][30]<= 127; ws[5][9 ][31]<=  23; ws[5][9 ][32]<= -57; ws[5][9 ][33]<=  15; ws[5][9 ][34]<= -17; ws[5][9 ][35]<= -72; ws[5][9 ][36]<= -73; ws[5][9 ][37]<=  38; ws[5][9 ][38]<= -16; ws[5][9 ][39]<=-150; ws[5][9 ][40]<=  22; ws[5][9 ][41]<=  48; ws[5][9 ][42]<=-227; ws[5][9 ][43]<= -88; ws[5][9 ][44]<=  29; ws[5][9 ][45]<=   4; ws[5][9 ][46]<=-204; ws[5][9 ][47]<=-110; ws[5][9 ][48]<= -61;
        ws[5][10][0]<=  73; ws[5][10][1]<= 151; ws[5][10][2]<= 115; ws[5][10][3]<= -89; ws[5][10][4]<=-127; ws[5][10][5]<=   0; ws[5][10][6]<=-105; ws[5][10][7]<= 145; ws[5][10][8]<=  18; ws[5][10][9]<=  -7; ws[5][10][10]<=-108; ws[5][10][11]<= -27; ws[5][10][12]<= 101; ws[5][10][13]<= -56; ws[5][10][14]<= 175; ws[5][10][15]<= -31; ws[5][10][16]<= -62; ws[5][10][17]<= -50; ws[5][10][18]<=  -5; ws[5][10][19]<=  96; ws[5][10][20]<= -44; ws[5][10][21]<= 174; ws[5][10][22]<=  92; ws[5][10][23]<= -56; ws[5][10][24]<=  26; ws[5][10][25]<=  20; ws[5][10][26]<=  22; ws[5][10][27]<= -57; ws[5][10][28]<= 194; ws[5][10][29]<= 154; ws[5][10][30]<=  30; ws[5][10][31]<=  18; ws[5][10][32]<= -16; ws[5][10][33]<=  -6; ws[5][10][34]<=  22; ws[5][10][35]<= 261; ws[5][10][36]<=  97; ws[5][10][37]<=  20; ws[5][10][38]<= -11; ws[5][10][39]<= -32; ws[5][10][40]<= -33; ws[5][10][41]<=  10; ws[5][10][42]<= 220; ws[5][10][43]<=  69; ws[5][10][44]<= -62; ws[5][10][45]<=-171; ws[5][10][46]<=-165; ws[5][10][47]<=  11; ws[5][10][48]<=  52;
        ws[5][11][0]<= 201; ws[5][11][1]<= 171; ws[5][11][2]<= 115; ws[5][11][3]<=  93; ws[5][11][4]<=  50; ws[5][11][5]<=  66; ws[5][11][6]<= 297; ws[5][11][7]<=  70; ws[5][11][8]<=  46; ws[5][11][9]<= -11; ws[5][11][10]<=  31; ws[5][11][11]<=  22; ws[5][11][12]<= -48; ws[5][11][13]<= 155; ws[5][11][14]<= 178; ws[5][11][15]<=   3; ws[5][11][16]<=  41; ws[5][11][17]<=  76; ws[5][11][18]<=  46; ws[5][11][19]<=  19; ws[5][11][20]<= 158; ws[5][11][21]<= 118; ws[5][11][22]<=  59; ws[5][11][23]<=  92; ws[5][11][24]<=  25; ws[5][11][25]<=  50; ws[5][11][26]<= -58; ws[5][11][27]<= 166; ws[5][11][28]<=  71; ws[5][11][29]<= 104; ws[5][11][30]<= 145; ws[5][11][31]<=  75; ws[5][11][32]<=  13; ws[5][11][33]<= -93; ws[5][11][34]<= 145; ws[5][11][35]<=   2; ws[5][11][36]<= -27; ws[5][11][37]<= 122; ws[5][11][38]<= 116; ws[5][11][39]<=   3; ws[5][11][40]<= -19; ws[5][11][41]<= 225; ws[5][11][42]<=-100; ws[5][11][43]<= -52; ws[5][11][44]<= 146; ws[5][11][45]<= 201; ws[5][11][46]<= 156; ws[5][11][47]<= 289; ws[5][11][48]<= 613;
        ws[5][12][0]<=  -4; ws[5][12][1]<=  19; ws[5][12][2]<= -21; ws[5][12][3]<=  47; ws[5][12][4]<=  14; ws[5][12][5]<= -46; ws[5][12][6]<=   9; ws[5][12][7]<=   0; ws[5][12][8]<=  -7; ws[5][12][9]<= -35; ws[5][12][10]<=  34; ws[5][12][11]<=   6; ws[5][12][12]<= -49; ws[5][12][13]<= -16; ws[5][12][14]<= -17; ws[5][12][15]<= -82; ws[5][12][16]<= -44; ws[5][12][17]<=  13; ws[5][12][18]<= -56; ws[5][12][19]<= -43; ws[5][12][20]<= -79; ws[5][12][21]<=-102; ws[5][12][22]<= -46; ws[5][12][23]<=  -8; ws[5][12][24]<=   9; ws[5][12][25]<= -48; ws[5][12][26]<=-110; ws[5][12][27]<=-101; ws[5][12][28]<= -53; ws[5][12][29]<=-114; ws[5][12][30]<= -58; ws[5][12][31]<= -12; ws[5][12][32]<= -47; ws[5][12][33]<=-109; ws[5][12][34]<=-154; ws[5][12][35]<=-100; ws[5][12][36]<= -55; ws[5][12][37]<= -33; ws[5][12][38]<= -42; ws[5][12][39]<= -11; ws[5][12][40]<=-158; ws[5][12][41]<=-191; ws[5][12][42]<= -70; ws[5][12][43]<= -74; ws[5][12][44]<=  -1; ws[5][12][45]<=  12; ws[5][12][46]<=  15; ws[5][12][47]<=-106; ws[5][12][48]<=-195;
        ws[5][13][0]<=  65; ws[5][13][1]<= 176; ws[5][13][2]<= 175; ws[5][13][3]<= 175; ws[5][13][4]<= 208; ws[5][13][5]<= 188; ws[5][13][6]<= 298; ws[5][13][7]<=  42; ws[5][13][8]<= 157; ws[5][13][9]<=  89; ws[5][13][10]<=  68; ws[5][13][11]<=   0; ws[5][13][12]<=  41; ws[5][13][13]<= 195; ws[5][13][14]<=  76; ws[5][13][15]<= 128; ws[5][13][16]<= 135; ws[5][13][17]<= -28; ws[5][13][18]<= -37; ws[5][13][19]<=  36; ws[5][13][20]<= 186; ws[5][13][21]<=  41; ws[5][13][22]<= 125; ws[5][13][23]<= 170; ws[5][13][24]<=  71; ws[5][13][25]<=-123; ws[5][13][26]<=   9; ws[5][13][27]<= 170; ws[5][13][28]<=  -6; ws[5][13][29]<=  -2; ws[5][13][30]<=  54; ws[5][13][31]<=  38; ws[5][13][32]<= -52; ws[5][13][33]<= -60; ws[5][13][34]<=  56; ws[5][13][35]<= -54; ws[5][13][36]<=  -3; ws[5][13][37]<= -27; ws[5][13][38]<=   5; ws[5][13][39]<= -57; ws[5][13][40]<= -40; ws[5][13][41]<=  19; ws[5][13][42]<=  52; ws[5][13][43]<=  32; ws[5][13][44]<=  26; ws[5][13][45]<= -14; ws[5][13][46]<=  23; ws[5][13][47]<= -60; ws[5][13][48]<= -81;
        ws[5][14][0]<=  49; ws[5][14][1]<=-102; ws[5][14][2]<=-163; ws[5][14][3]<= -25; ws[5][14][4]<= 134; ws[5][14][5]<=  91; ws[5][14][6]<= 223; ws[5][14][7]<=  17; ws[5][14][8]<=-174; ws[5][14][9]<= -92; ws[5][14][10]<=  39; ws[5][14][11]<= 111; ws[5][14][12]<= 111; ws[5][14][13]<= 105; ws[5][14][14]<=  10; ws[5][14][15]<= -71; ws[5][14][16]<= -72; ws[5][14][17]<=  68; ws[5][14][18]<= 111; ws[5][14][19]<=  99; ws[5][14][20]<=  80; ws[5][14][21]<=  54; ws[5][14][22]<=  78; ws[5][14][23]<=  76; ws[5][14][24]<=  65; ws[5][14][25]<=  23; ws[5][14][26]<=  97; ws[5][14][27]<= 128; ws[5][14][28]<= 157; ws[5][14][29]<= 174; ws[5][14][30]<=  42; ws[5][14][31]<=  44; ws[5][14][32]<= -54; ws[5][14][33]<=  11; ws[5][14][34]<= 179; ws[5][14][35]<=  11; ws[5][14][36]<= 174; ws[5][14][37]<=  90; ws[5][14][38]<= -16; ws[5][14][39]<=-126; ws[5][14][40]<= -25; ws[5][14][41]<= 229; ws[5][14][42]<= -71; ws[5][14][43]<=  26; ws[5][14][44]<= 113; ws[5][14][45]<=-129; ws[5][14][46]<=-205; ws[5][14][47]<=-148; ws[5][14][48]<=  76;
        ws[5][15][0]<=  22; ws[5][15][1]<=  41; ws[5][15][2]<=  72; ws[5][15][3]<= 119; ws[5][15][4]<= 102; ws[5][15][5]<=  40; ws[5][15][6]<=  29; ws[5][15][7]<=   4; ws[5][15][8]<=  60; ws[5][15][9]<= 130; ws[5][15][10]<= 199; ws[5][15][11]<= 133; ws[5][15][12]<=  75; ws[5][15][13]<=  65; ws[5][15][14]<=  -8; ws[5][15][15]<=  40; ws[5][15][16]<= 126; ws[5][15][17]<= 157; ws[5][15][18]<= 149; ws[5][15][19]<=  71; ws[5][15][20]<=  62; ws[5][15][21]<= -23; ws[5][15][22]<= -24; ws[5][15][23]<=  84; ws[5][15][24]<=  61; ws[5][15][25]<=  70; ws[5][15][26]<= -12; ws[5][15][27]<= 106; ws[5][15][28]<=  39; ws[5][15][29]<=   7; ws[5][15][30]<= -29; ws[5][15][31]<=  28; ws[5][15][32]<=  47; ws[5][15][33]<=   3; ws[5][15][34]<=  72; ws[5][15][35]<= 119; ws[5][15][36]<=  -7; ws[5][15][37]<= -30; ws[5][15][38]<= -75; ws[5][15][39]<=  13; ws[5][15][40]<=  -3; ws[5][15][41]<= 158; ws[5][15][42]<= 164; ws[5][15][43]<= 135; ws[5][15][44]<=  14; ws[5][15][45]<= -96; ws[5][15][46]<=  22; ws[5][15][47]<=  59; ws[5][15][48]<= 186;

        ws[6][0 ][0]<= -58; ws[6][0 ][1]<= -87; ws[6][0 ][2]<= -73; ws[6][0 ][3]<=  18; ws[6][0 ][4]<= -76; ws[6][0 ][5]<=-145; ws[6][0 ][6]<=-187; ws[6][0 ][7]<= -49; ws[6][0 ][8]<= -44; ws[6][0 ][9]<= -49; ws[6][0 ][10]<=   0; ws[6][0 ][11]<= -28; ws[6][0 ][12]<=-115; ws[6][0 ][13]<=-130; ws[6][0 ][14]<= -40; ws[6][0 ][15]<= -54; ws[6][0 ][16]<= -31; ws[6][0 ][17]<= -28; ws[6][0 ][18]<= -32; ws[6][0 ][19]<= -72; ws[6][0 ][20]<=-103; ws[6][0 ][21]<= -79; ws[6][0 ][22]<= -25; ws[6][0 ][23]<= -60; ws[6][0 ][24]<= -55; ws[6][0 ][25]<= -66; ws[6][0 ][26]<= -92; ws[6][0 ][27]<= -59; ws[6][0 ][28]<=   7; ws[6][0 ][29]<= -77; ws[6][0 ][30]<= -72; ws[6][0 ][31]<= -36; ws[6][0 ][32]<=-110; ws[6][0 ][33]<= -84; ws[6][0 ][34]<=  -9; ws[6][0 ][35]<=  -5; ws[6][0 ][36]<= -22; ws[6][0 ][37]<= -65; ws[6][0 ][38]<=-132; ws[6][0 ][39]<=-100; ws[6][0 ][40]<= -41; ws[6][0 ][41]<=  -4; ws[6][0 ][42]<= -40; ws[6][0 ][43]<= -69; ws[6][0 ][44]<= -55; ws[6][0 ][45]<=-138; ws[6][0 ][46]<=-178; ws[6][0 ][47]<= -91; ws[6][0 ][48]<= -29;
        ws[6][1 ][0]<=-136; ws[6][1 ][1]<= -76; ws[6][1 ][2]<= -27; ws[6][1 ][3]<=  44; ws[6][1 ][4]<=  -4; ws[6][1 ][5]<= -58; ws[6][1 ][6]<=-151; ws[6][1 ][7]<= -60; ws[6][1 ][8]<= -58; ws[6][1 ][9]<= -10; ws[6][1 ][10]<= -81; ws[6][1 ][11]<= -59; ws[6][1 ][12]<= -54; ws[6][1 ][13]<=-105; ws[6][1 ][14]<= -33; ws[6][1 ][15]<=   6; ws[6][1 ][16]<=  49; ws[6][1 ][17]<=  32; ws[6][1 ][18]<=  -1; ws[6][1 ][19]<=  -5; ws[6][1 ][20]<= -26; ws[6][1 ][21]<= -19; ws[6][1 ][22]<=  20; ws[6][1 ][23]<=  36; ws[6][1 ][24]<=  31; ws[6][1 ][25]<=  54; ws[6][1 ][26]<=  81; ws[6][1 ][27]<= -29; ws[6][1 ][28]<= -12; ws[6][1 ][29]<=   6; ws[6][1 ][30]<=  24; ws[6][1 ][31]<= -48; ws[6][1 ][32]<=  35; ws[6][1 ][33]<=  35; ws[6][1 ][34]<=-123; ws[6][1 ][35]<= -26; ws[6][1 ][36]<=  18; ws[6][1 ][37]<= -38; ws[6][1 ][38]<= -80; ws[6][1 ][39]<=-102; ws[6][1 ][40]<=-112; ws[6][1 ][41]<=-216; ws[6][1 ][42]<=  39; ws[6][1 ][43]<= -25; ws[6][1 ][44]<= -67; ws[6][1 ][45]<=-145; ws[6][1 ][46]<=-191; ws[6][1 ][47]<=-202; ws[6][1 ][48]<=-248;
        ws[6][2 ][0]<=  45; ws[6][2 ][1]<=  32; ws[6][2 ][2]<=   1; ws[6][2 ][3]<= -48; ws[6][2 ][4]<= -50; ws[6][2 ][5]<= -43; ws[6][2 ][6]<=-220; ws[6][2 ][7]<= -11; ws[6][2 ][8]<=  -4; ws[6][2 ][9]<= -57; ws[6][2 ][10]<= -30; ws[6][2 ][11]<=  34; ws[6][2 ][12]<= 100; ws[6][2 ][13]<= -39; ws[6][2 ][14]<= -81; ws[6][2 ][15]<= -35; ws[6][2 ][16]<=-144; ws[6][2 ][17]<= -71; ws[6][2 ][18]<=  17; ws[6][2 ][19]<=  70; ws[6][2 ][20]<=  12; ws[6][2 ][21]<=-119; ws[6][2 ][22]<= -53; ws[6][2 ][23]<=-141; ws[6][2 ][24]<=-124; ws[6][2 ][25]<=  28; ws[6][2 ][26]<=  33; ws[6][2 ][27]<=   0; ws[6][2 ][28]<= -39; ws[6][2 ][29]<= -92; ws[6][2 ][30]<=-133; ws[6][2 ][31]<=-114; ws[6][2 ][32]<=  -5; ws[6][2 ][33]<=  19; ws[6][2 ][34]<=  52; ws[6][2 ][35]<= -66; ws[6][2 ][36]<= -66; ws[6][2 ][37]<=-106; ws[6][2 ][38]<=  -8; ws[6][2 ][39]<= 114; ws[6][2 ][40]<=  29; ws[6][2 ][41]<= -13; ws[6][2 ][42]<= -30; ws[6][2 ][43]<=-137; ws[6][2 ][44]<= -97; ws[6][2 ][45]<=  21; ws[6][2 ][46]<=  52; ws[6][2 ][47]<= -31; ws[6][2 ][48]<= -80;
        ws[6][3 ][0]<= -11; ws[6][3 ][1]<= -75; ws[6][3 ][2]<= -99; ws[6][3 ][3]<= -83; ws[6][3 ][4]<= -64; ws[6][3 ][5]<= -28; ws[6][3 ][6]<=  34; ws[6][3 ][7]<= -43; ws[6][3 ][8]<=  11; ws[6][3 ][9]<=  61; ws[6][3 ][10]<=  52; ws[6][3 ][11]<= -38; ws[6][3 ][12]<= -79; ws[6][3 ][13]<=  75; ws[6][3 ][14]<=  45; ws[6][3 ][15]<= -14; ws[6][3 ][16]<= 136; ws[6][3 ][17]<= 122; ws[6][3 ][18]<= -21; ws[6][3 ][19]<=-134; ws[6][3 ][20]<=  28; ws[6][3 ][21]<= 212; ws[6][3 ][22]<=  88; ws[6][3 ][23]<= 181; ws[6][3 ][24]<= 136; ws[6][3 ][25]<=  10; ws[6][3 ][26]<=-131; ws[6][3 ][27]<=  90; ws[6][3 ][28]<= 344; ws[6][3 ][29]<=  92; ws[6][3 ][30]<= 161; ws[6][3 ][31]<=   3; ws[6][3 ][32]<=  -2; ws[6][3 ][33]<= -86; ws[6][3 ][34]<= 152; ws[6][3 ][35]<= 155; ws[6][3 ][36]<=   3; ws[6][3 ][37]<=  20; ws[6][3 ][38]<=  -6; ws[6][3 ][39]<= -36; ws[6][3 ][40]<=  15; ws[6][3 ][41]<= 181; ws[6][3 ][42]<=  10; ws[6][3 ][43]<= -82; ws[6][3 ][44]<= -45; ws[6][3 ][45]<=-220; ws[6][3 ][46]<=-100; ws[6][3 ][47]<= -18; ws[6][3 ][48]<=  51;
        ws[6][4 ][0]<=  74; ws[6][4 ][1]<=   5; ws[6][4 ][2]<= -61; ws[6][4 ][3]<=-101; ws[6][4 ][4]<= -36; ws[6][4 ][5]<=  43; ws[6][4 ][6]<=-287; ws[6][4 ][7]<=   0; ws[6][4 ][8]<=  -7; ws[6][4 ][9]<= -27; ws[6][4 ][10]<= -41; ws[6][4 ][11]<= -23; ws[6][4 ][12]<=  62; ws[6][4 ][13]<=-147; ws[6][4 ][14]<= -65; ws[6][4 ][15]<=   1; ws[6][4 ][16]<= -77; ws[6][4 ][17]<=  62; ws[6][4 ][18]<=  34; ws[6][4 ][19]<=  47; ws[6][4 ][20]<=-108; ws[6][4 ][21]<=   0; ws[6][4 ][22]<= -15; ws[6][4 ][23]<=-117; ws[6][4 ][24]<= -55; ws[6][4 ][25]<=  -4; ws[6][4 ][26]<=  25; ws[6][4 ][27]<=-110; ws[6][4 ][28]<=   9; ws[6][4 ][29]<= 101; ws[6][4 ][30]<=-130; ws[6][4 ][31]<=-133; ws[6][4 ][32]<= -66; ws[6][4 ][33]<= -51; ws[6][4 ][34]<=-108; ws[6][4 ][35]<= -11; ws[6][4 ][36]<=  87; ws[6][4 ][37]<= -83; ws[6][4 ][38]<=-129; ws[6][4 ][39]<=-137; ws[6][4 ][40]<=-109; ws[6][4 ][41]<=-100; ws[6][4 ][42]<= -26; ws[6][4 ][43]<=  67; ws[6][4 ][44]<= -33; ws[6][4 ][45]<= -82; ws[6][4 ][46]<=-169; ws[6][4 ][47]<=-146; ws[6][4 ][48]<= -82;
        ws[6][5 ][0]<=-134; ws[6][5 ][1]<= -48; ws[6][5 ][2]<= -54; ws[6][5 ][3]<= -61; ws[6][5 ][4]<=-172; ws[6][5 ][5]<= -33; ws[6][5 ][6]<=  37; ws[6][5 ][7]<=-122; ws[6][5 ][8]<= -87; ws[6][5 ][9]<= -30; ws[6][5 ][10]<= -65; ws[6][5 ][11]<=-192; ws[6][5 ][12]<= -44; ws[6][5 ][13]<=  72; ws[6][5 ][14]<= -36; ws[6][5 ][15]<= -69; ws[6][5 ][16]<= -15; ws[6][5 ][17]<= -34; ws[6][5 ][18]<=-201; ws[6][5 ][19]<=  -2; ws[6][5 ][20]<=  62; ws[6][5 ][21]<=   0; ws[6][5 ][22]<= -44; ws[6][5 ][23]<= -11; ws[6][5 ][24]<= -35; ws[6][5 ][25]<=-214; ws[6][5 ][26]<= -76; ws[6][5 ][27]<=  19; ws[6][5 ][28]<=  93; ws[6][5 ][29]<= -43; ws[6][5 ][30]<=  36; ws[6][5 ][31]<=  48; ws[6][5 ][32]<=-153; ws[6][5 ][33]<=-143; ws[6][5 ][34]<=  70; ws[6][5 ][35]<= 135; ws[6][5 ][36]<=  23; ws[6][5 ][37]<= -21; ws[6][5 ][38]<=  62; ws[6][5 ][39]<= -87; ws[6][5 ][40]<=-105; ws[6][5 ][41]<= 163; ws[6][5 ][42]<=  45; ws[6][5 ][43]<= -38; ws[6][5 ][44]<= -39; ws[6][5 ][45]<=  37; ws[6][5 ][46]<= -70; ws[6][5 ][47]<=-118; ws[6][5 ][48]<= 123;
        ws[6][6 ][0]<= 124; ws[6][6 ][1]<=  44; ws[6][6 ][2]<=  26; ws[6][6 ][3]<= 105; ws[6][6 ][4]<= 168; ws[6][6 ][5]<=  63; ws[6][6 ][6]<=-130; ws[6][6 ][7]<= -36; ws[6][6 ][8]<= -39; ws[6][6 ][9]<= -40; ws[6][6 ][10]<= -97; ws[6][6 ][11]<= 109; ws[6][6 ][12]<=  30; ws[6][6 ][13]<= -71; ws[6][6 ][14]<=-166; ws[6][6 ][15]<= -73; ws[6][6 ][16]<=-128; ws[6][6 ][17]<=-107; ws[6][6 ][18]<=  50; ws[6][6 ][19]<= 125; ws[6][6 ][20]<=   2; ws[6][6 ][21]<=-166; ws[6][6 ][22]<= -63; ws[6][6 ][23]<= -68; ws[6][6 ][24]<= -49; ws[6][6 ][25]<=  -8; ws[6][6 ][26]<= 134; ws[6][6 ][27]<=  71; ws[6][6 ][28]<=-230; ws[6][6 ][29]<= -32; ws[6][6 ][30]<=  25; ws[6][6 ][31]<=  16; ws[6][6 ][32]<=-138; ws[6][6 ][33]<= -16; ws[6][6 ][34]<= -13; ws[6][6 ][35]<=-112; ws[6][6 ][36]<=  -8; ws[6][6 ][37]<=  59; ws[6][6 ][38]<=  78; ws[6][6 ][39]<=-167; ws[6][6 ][40]<=-142; ws[6][6 ][41]<= -80; ws[6][6 ][42]<=  98; ws[6][6 ][43]<=  73; ws[6][6 ][44]<=   2; ws[6][6 ][45]<=  34; ws[6][6 ][46]<=-182; ws[6][6 ][47]<=-244; ws[6][6 ][48]<= -68;
        ws[6][7 ][0]<= 136; ws[6][7 ][1]<=   4; ws[6][7 ][2]<=  20; ws[6][7 ][3]<=  43; ws[6][7 ][4]<= -74; ws[6][7 ][5]<=   0; ws[6][7 ][6]<= 183; ws[6][7 ][7]<= 101; ws[6][7 ][8]<= -31; ws[6][7 ][9]<=  12; ws[6][7 ][10]<=  59; ws[6][7 ][11]<= -49; ws[6][7 ][12]<= -26; ws[6][7 ][13]<= 165; ws[6][7 ][14]<=  76; ws[6][7 ][15]<= -36; ws[6][7 ][16]<=   0; ws[6][7 ][17]<=  52; ws[6][7 ][18]<=  11; ws[6][7 ][19]<= -39; ws[6][7 ][20]<=  26; ws[6][7 ][21]<=  47; ws[6][7 ][22]<= -26; ws[6][7 ][23]<=-125; ws[6][7 ][24]<= -61; ws[6][7 ][25]<= -76; ws[6][7 ][26]<=-109; ws[6][7 ][27]<=-150; ws[6][7 ][28]<= 165; ws[6][7 ][29]<=  61; ws[6][7 ][30]<= -34; ws[6][7 ][31]<=  39; ws[6][7 ][32]<=  63; ws[6][7 ][33]<=   3; ws[6][7 ][34]<=-163; ws[6][7 ][35]<= 165; ws[6][7 ][36]<=  38; ws[6][7 ][37]<= -99; ws[6][7 ][38]<=  24; ws[6][7 ][39]<=  43; ws[6][7 ][40]<= -24; ws[6][7 ][41]<=-190; ws[6][7 ][42]<= 112; ws[6][7 ][43]<= -42; ws[6][7 ][44]<=-169; ws[6][7 ][45]<=-161; ws[6][7 ][46]<=-183; ws[6][7 ][47]<=-208; ws[6][7 ][48]<=-159;
        ws[6][8 ][0]<=   5; ws[6][8 ][1]<=  62; ws[6][8 ][2]<= 113; ws[6][8 ][3]<=  57; ws[6][8 ][4]<=  49; ws[6][8 ][5]<= 116; ws[6][8 ][6]<=  18; ws[6][8 ][7]<=   0; ws[6][8 ][8]<=  65; ws[6][8 ][9]<= 114; ws[6][8 ][10]<=  11; ws[6][8 ][11]<=-102; ws[6][8 ][12]<= -35; ws[6][8 ][13]<= -34; ws[6][8 ][14]<= -15; ws[6][8 ][15]<=  64; ws[6][8 ][16]<=  60; ws[6][8 ][17]<= -61; ws[6][8 ][18]<=-217; ws[6][8 ][19]<=-126; ws[6][8 ][20]<= -14; ws[6][8 ][21]<= -35; ws[6][8 ][22]<= -64; ws[6][8 ][23]<= -22; ws[6][8 ][24]<=-179; ws[6][8 ][25]<=-222; ws[6][8 ][26]<=-181; ws[6][8 ][27]<= -15; ws[6][8 ][28]<= -47; ws[6][8 ][29]<= -70; ws[6][8 ][30]<=  10; ws[6][8 ][31]<=-151; ws[6][8 ][32]<=-214; ws[6][8 ][33]<=-128; ws[6][8 ][34]<=  -2; ws[6][8 ][35]<=  87; ws[6][8 ][36]<= -20; ws[6][8 ][37]<= -10; ws[6][8 ][38]<=-105; ws[6][8 ][39]<=-177; ws[6][8 ][40]<=-129; ws[6][8 ][41]<=  -1; ws[6][8 ][42]<= 300; ws[6][8 ][43]<= 125; ws[6][8 ][44]<= 168; ws[6][8 ][45]<= -48; ws[6][8 ][46]<=-153; ws[6][8 ][47]<=-272; ws[6][8 ][48]<=  13;
        ws[6][9 ][0]<=-136; ws[6][9 ][1]<=-134; ws[6][9 ][2]<=-206; ws[6][9 ][3]<=-179; ws[6][9 ][4]<=-119; ws[6][9 ][5]<=  10; ws[6][9 ][6]<=  -6; ws[6][9 ][7]<= -63; ws[6][9 ][8]<= -35; ws[6][9 ][9]<= -53; ws[6][9 ][10]<= -99; ws[6][9 ][11]<= -49; ws[6][9 ][12]<=  51; ws[6][9 ][13]<= 128; ws[6][9 ][14]<= -15; ws[6][9 ][15]<=  44; ws[6][9 ][16]<=  19; ws[6][9 ][17]<= -41; ws[6][9 ][18]<=  60; ws[6][9 ][19]<= 122; ws[6][9 ][20]<= 147; ws[6][9 ][21]<= -12; ws[6][9 ][22]<=  12; ws[6][9 ][23]<=  -5; ws[6][9 ][24]<=  11; ws[6][9 ][25]<=  61; ws[6][9 ][26]<=  63; ws[6][9 ][27]<= 167; ws[6][9 ][28]<= -60; ws[6][9 ][29]<=  12; ws[6][9 ][30]<= -13; ws[6][9 ][31]<=   9; ws[6][9 ][32]<=  80; ws[6][9 ][33]<=  50; ws[6][9 ][34]<= 130; ws[6][9 ][35]<= -80; ws[6][9 ][36]<= -57; ws[6][9 ][37]<=  -1; ws[6][9 ][38]<= -13; ws[6][9 ][39]<=   1; ws[6][9 ][40]<= -50; ws[6][9 ][41]<=  26; ws[6][9 ][42]<=-226; ws[6][9 ][43]<=-198; ws[6][9 ][44]<=-118; ws[6][9 ][45]<= -68; ws[6][9 ][46]<= -98; ws[6][9 ][47]<= -83; ws[6][9 ][48]<=-120;
        ws[6][10][0]<=-110; ws[6][10][1]<= -24; ws[6][10][2]<= -41; ws[6][10][3]<=  17; ws[6][10][4]<=  21; ws[6][10][5]<= -79; ws[6][10][6]<=-288; ws[6][10][7]<= -66; ws[6][10][8]<=  13; ws[6][10][9]<=  15; ws[6][10][10]<=   4; ws[6][10][11]<=  49; ws[6][10][12]<= -65; ws[6][10][13]<=-175; ws[6][10][14]<=  26; ws[6][10][15]<= 143; ws[6][10][16]<=  91; ws[6][10][17]<=  -8; ws[6][10][18]<=   8; ws[6][10][19]<= -35; ws[6][10][20]<=-159; ws[6][10][21]<=  52; ws[6][10][22]<=  96; ws[6][10][23]<=  55; ws[6][10][24]<= -32; ws[6][10][25]<=  10; ws[6][10][26]<=   6; ws[6][10][27]<=-119; ws[6][10][28]<=  43; ws[6][10][29]<=  88; ws[6][10][30]<= 106; ws[6][10][31]<= -17; ws[6][10][32]<=   8; ws[6][10][33]<= -49; ws[6][10][34]<=-160; ws[6][10][35]<= 100; ws[6][10][36]<= 114; ws[6][10][37]<= 139; ws[6][10][38]<= -26; ws[6][10][39]<= -46; ws[6][10][40]<= -92; ws[6][10][41]<=-128; ws[6][10][42]<= 106; ws[6][10][43]<=  97; ws[6][10][44]<= 146; ws[6][10][45]<=   6; ws[6][10][46]<=-120; ws[6][10][47]<=-159; ws[6][10][48]<=-107;
        ws[6][11][0]<= -98; ws[6][11][1]<= -41; ws[6][11][2]<=-144; ws[6][11][3]<=-131; ws[6][11][4]<= -14; ws[6][11][5]<=  51; ws[6][11][6]<= 105; ws[6][11][7]<= -38; ws[6][11][8]<=  53; ws[6][11][9]<=-133; ws[6][11][10]<=-163; ws[6][11][11]<= -80; ws[6][11][12]<=  54; ws[6][11][13]<= 126; ws[6][11][14]<=-114; ws[6][11][15]<=  16; ws[6][11][16]<=-149; ws[6][11][17]<=-190; ws[6][11][18]<= -79; ws[6][11][19]<= -21; ws[6][11][20]<=  88; ws[6][11][21]<= -43; ws[6][11][22]<=  49; ws[6][11][23]<= -52; ws[6][11][24]<=-104; ws[6][11][25]<=  -7; ws[6][11][26]<= 105; ws[6][11][27]<=  77; ws[6][11][28]<= -30; ws[6][11][29]<=  68; ws[6][11][30]<= -16; ws[6][11][31]<= -23; ws[6][11][32]<=   7; ws[6][11][33]<=  72; ws[6][11][34]<=  90; ws[6][11][35]<=   1; ws[6][11][36]<=   3; ws[6][11][37]<= -60; ws[6][11][38]<= -55; ws[6][11][39]<=  47; ws[6][11][40]<=  87; ws[6][11][41]<=  63; ws[6][11][42]<= -33; ws[6][11][43]<= -83; ws[6][11][44]<=-180; ws[6][11][45]<= -44; ws[6][11][46]<=  80; ws[6][11][47]<= -34; ws[6][11][48]<=  19;
        ws[6][12][0]<= -87; ws[6][12][1]<=  15; ws[6][12][2]<=  -9; ws[6][12][3]<= 104; ws[6][12][4]<= 163; ws[6][12][5]<=  32; ws[6][12][6]<=  -9; ws[6][12][7]<= -73; ws[6][12][8]<=  -1; ws[6][12][9]<= -12; ws[6][12][10]<=  33; ws[6][12][11]<=  52; ws[6][12][12]<=  31; ws[6][12][13]<=  14; ws[6][12][14]<= -65; ws[6][12][15]<= -62; ws[6][12][16]<=-109; ws[6][12][17]<=-111; ws[6][12][18]<= -48; ws[6][12][19]<=  13; ws[6][12][20]<=  13; ws[6][12][21]<= -99; ws[6][12][22]<= -80; ws[6][12][23]<= -69; ws[6][12][24]<=-176; ws[6][12][25]<= -32; ws[6][12][26]<=  -5; ws[6][12][27]<= -56; ws[6][12][28]<=-109; ws[6][12][29]<=  -7; ws[6][12][30]<= -87; ws[6][12][31]<=-220; ws[6][12][32]<= -80; ws[6][12][33]<= -57; ws[6][12][34]<=-151; ws[6][12][35]<=-128; ws[6][12][36]<= -23; ws[6][12][37]<= -64; ws[6][12][38]<=-134; ws[6][12][39]<= -92; ws[6][12][40]<= -83; ws[6][12][41]<=-177; ws[6][12][42]<=-135; ws[6][12][43]<=  33; ws[6][12][44]<= -53; ws[6][12][45]<= -77; ws[6][12][46]<=-101; ws[6][12][47]<= -93; ws[6][12][48]<=-132;
        ws[6][13][0]<= 169; ws[6][13][1]<= 116; ws[6][13][2]<= 126; ws[6][13][3]<= 131; ws[6][13][4]<=  72; ws[6][13][5]<=  89; ws[6][13][6]<=  51; ws[6][13][7]<=  96; ws[6][13][8]<= 126; ws[6][13][9]<= 114; ws[6][13][10]<=  67; ws[6][13][11]<=  41; ws[6][13][12]<=  59; ws[6][13][13]<= -61; ws[6][13][14]<= 108; ws[6][13][15]<=  75; ws[6][13][16]<= 142; ws[6][13][17]<=  41; ws[6][13][18]<=  87; ws[6][13][19]<=   3; ws[6][13][20]<= -19; ws[6][13][21]<= 104; ws[6][13][22]<=  45; ws[6][13][23]<=  62; ws[6][13][24]<=  24; ws[6][13][25]<=  48; ws[6][13][26]<=   0; ws[6][13][27]<= -46; ws[6][13][28]<=  82; ws[6][13][29]<= -42; ws[6][13][30]<= -35; ws[6][13][31]<=  13; ws[6][13][32]<=  48; ws[6][13][33]<=  38; ws[6][13][34]<= -78; ws[6][13][35]<=  69; ws[6][13][36]<=   7; ws[6][13][37]<= -39; ws[6][13][38]<= -20; ws[6][13][39]<=  64; ws[6][13][40]<=  19; ws[6][13][41]<= -21; ws[6][13][42]<= 223; ws[6][13][43]<= 134; ws[6][13][44]<= 110; ws[6][13][45]<=  67; ws[6][13][46]<= 132; ws[6][13][47]<=  59; ws[6][13][48]<= -53;
        ws[6][14][0]<=-221; ws[6][14][1]<=-147; ws[6][14][2]<=-174; ws[6][14][3]<=-174; ws[6][14][4]<=-140; ws[6][14][5]<=-195; ws[6][14][6]<=-239; ws[6][14][7]<=   3; ws[6][14][8]<=  63; ws[6][14][9]<=  86; ws[6][14][10]<=  50; ws[6][14][11]<=  39; ws[6][14][12]<= -33; ws[6][14][13]<=-173; ws[6][14][14]<= -13; ws[6][14][15]<=  59; ws[6][14][16]<=  57; ws[6][14][17]<= -12; ws[6][14][18]<=  36; ws[6][14][19]<=  29; ws[6][14][20]<=-183; ws[6][14][21]<= -53; ws[6][14][22]<=   1; ws[6][14][23]<=   3; ws[6][14][24]<= -85; ws[6][14][25]<=  -5; ws[6][14][26]<= -34; ws[6][14][27]<=-141; ws[6][14][28]<= -49; ws[6][14][29]<=  53; ws[6][14][30]<=  22; ws[6][14][31]<=  -3; ws[6][14][32]<=  23; ws[6][14][33]<=  61; ws[6][14][34]<=-137; ws[6][14][35]<= -88; ws[6][14][36]<=  17; ws[6][14][37]<=  63; ws[6][14][38]<=  43; ws[6][14][39]<=  25; ws[6][14][40]<=  -3; ws[6][14][41]<=-110; ws[6][14][42]<=-342; ws[6][14][43]<=-133; ws[6][14][44]<= -69; ws[6][14][45]<=-108; ws[6][14][46]<=-117; ws[6][14][47]<=-137; ws[6][14][48]<=-274;
        ws[6][15][0]<=  58; ws[6][15][1]<= 124; ws[6][15][2]<= -19; ws[6][15][3]<= -49; ws[6][15][4]<= -72; ws[6][15][5]<=-119; ws[6][15][6]<=-184; ws[6][15][7]<=  15; ws[6][15][8]<=  90; ws[6][15][9]<= -25; ws[6][15][10]<= -37; ws[6][15][11]<= -72; ws[6][15][12]<=-123; ws[6][15][13]<= -74; ws[6][15][14]<=  67; ws[6][15][15]<=  78; ws[6][15][16]<= -89; ws[6][15][17]<=  26; ws[6][15][18]<= -35; ws[6][15][19]<=-172; ws[6][15][20]<=  19; ws[6][15][21]<= -10; ws[6][15][22]<=  55; ws[6][15][23]<= -75; ws[6][15][24]<= -38; ws[6][15][25]<=-159; ws[6][15][26]<=-199; ws[6][15][27]<=  33; ws[6][15][28]<=  43; ws[6][15][29]<=  30; ws[6][15][30]<= -81; ws[6][15][31]<=-100; ws[6][15][32]<=-103; ws[6][15][33]<=-104; ws[6][15][34]<=  49; ws[6][15][35]<=  -3; ws[6][15][36]<= -27; ws[6][15][37]<= -80; ws[6][15][38]<= -29; ws[6][15][39]<= -45; ws[6][15][40]<=  12; ws[6][15][41]<= 161; ws[6][15][42]<=  99; ws[6][15][43]<=  40; ws[6][15][44]<=  -2; ws[6][15][45]<=  41; ws[6][15][46]<=  78; ws[6][15][47]<= 190; ws[6][15][48]<= 314;

        ws[7][0 ][0]<= -29; ws[7][0 ][1]<=  44; ws[7][0 ][2]<=  27; ws[7][0 ][3]<= -92; ws[7][0 ][4]<=  -8; ws[7][0 ][5]<= -81; ws[7][0 ][6]<= -13; ws[7][0 ][7]<=-184; ws[7][0 ][8]<=  42; ws[7][0 ][9]<=  20; ws[7][0 ][10]<=-100; ws[7][0 ][11]<=   8; ws[7][0 ][12]<=   8; ws[7][0 ][13]<=   6; ws[7][0 ][14]<=  15; ws[7][0 ][15]<=  -9; ws[7][0 ][16]<= -45; ws[7][0 ][17]<= -67; ws[7][0 ][18]<= -17; ws[7][0 ][19]<= -12; ws[7][0 ][20]<= -69; ws[7][0 ][21]<= -44; ws[7][0 ][22]<= -78; ws[7][0 ][23]<= -43; ws[7][0 ][24]<= -44; ws[7][0 ][25]<= -64; ws[7][0 ][26]<= -55; ws[7][0 ][27]<=-145; ws[7][0 ][28]<= -72; ws[7][0 ][29]<= -33; ws[7][0 ][30]<= -81; ws[7][0 ][31]<= -17; ws[7][0 ][32]<=-141; ws[7][0 ][33]<= -52; ws[7][0 ][34]<= -86; ws[7][0 ][35]<= -78; ws[7][0 ][36]<= -48; ws[7][0 ][37]<= -54; ws[7][0 ][38]<= -87; ws[7][0 ][39]<=-136; ws[7][0 ][40]<=  12; ws[7][0 ][41]<= -14; ws[7][0 ][42]<=-114; ws[7][0 ][43]<= -23; ws[7][0 ][44]<=-110; ws[7][0 ][45]<= -40; ws[7][0 ][46]<= -86; ws[7][0 ][47]<= -42; ws[7][0 ][48]<= -16;
        ws[7][1 ][0]<=  11; ws[7][1 ][1]<=  79; ws[7][1 ][2]<= -14; ws[7][1 ][3]<=  43; ws[7][1 ][4]<=   4; ws[7][1 ][5]<= -79; ws[7][1 ][6]<= -79; ws[7][1 ][7]<=-103; ws[7][1 ][8]<= 108; ws[7][1 ][9]<= 230; ws[7][1 ][10]<=  45; ws[7][1 ][11]<=  24; ws[7][1 ][12]<= -75; ws[7][1 ][13]<=  11; ws[7][1 ][14]<= -78; ws[7][1 ][15]<=   1; ws[7][1 ][16]<= 220; ws[7][1 ][17]<= 111; ws[7][1 ][18]<=  18; ws[7][1 ][19]<= -49; ws[7][1 ][20]<=  51; ws[7][1 ][21]<= -48; ws[7][1 ][22]<=  78; ws[7][1 ][23]<= 181; ws[7][1 ][24]<= 206; ws[7][1 ][25]<=  33; ws[7][1 ][26]<=  11; ws[7][1 ][27]<=  94; ws[7][1 ][28]<=  44; ws[7][1 ][29]<=  32; ws[7][1 ][30]<=  81; ws[7][1 ][31]<= 157; ws[7][1 ][32]<=  13; ws[7][1 ][33]<= -27; ws[7][1 ][34]<= -23; ws[7][1 ][35]<=  69; ws[7][1 ][36]<= -21; ws[7][1 ][37]<= -75; ws[7][1 ][38]<= 107; ws[7][1 ][39]<=  55; ws[7][1 ][40]<= -25; ws[7][1 ][41]<= -15; ws[7][1 ][42]<= 156; ws[7][1 ][43]<=-147; ws[7][1 ][44]<=-264; ws[7][1 ][45]<=  37; ws[7][1 ][46]<=  50; ws[7][1 ][47]<= -29; ws[7][1 ][48]<= -13;
        ws[7][2 ][0]<= -48; ws[7][2 ][1]<= -26; ws[7][2 ][2]<=-110; ws[7][2 ][3]<=-109; ws[7][2 ][4]<= -64; ws[7][2 ][5]<=  22; ws[7][2 ][6]<=  57; ws[7][2 ][7]<=-108; ws[7][2 ][8]<= -44; ws[7][2 ][9]<= -90; ws[7][2 ][10]<= -31; ws[7][2 ][11]<= -38; ws[7][2 ][12]<= -69; ws[7][2 ][13]<=  42; ws[7][2 ][14]<= -39; ws[7][2 ][15]<= -95; ws[7][2 ][16]<=-125; ws[7][2 ][17]<=   8; ws[7][2 ][18]<=  18; ws[7][2 ][19]<= -29; ws[7][2 ][20]<= -25; ws[7][2 ][21]<=   4; ws[7][2 ][22]<= -78; ws[7][2 ][23]<= -70; ws[7][2 ][24]<=  -9; ws[7][2 ][25]<=   8; ws[7][2 ][26]<= -96; ws[7][2 ][27]<= -47; ws[7][2 ][28]<= -53; ws[7][2 ][29]<= -61; ws[7][2 ][30]<= -99; ws[7][2 ][31]<=  26; ws[7][2 ][32]<=  20; ws[7][2 ][33]<= -68; ws[7][2 ][34]<= -81; ws[7][2 ][35]<= -87; ws[7][2 ][36]<= -47; ws[7][2 ][37]<= -82; ws[7][2 ][38]<= -25; ws[7][2 ][39]<= -83; ws[7][2 ][40]<= -73; ws[7][2 ][41]<= -27; ws[7][2 ][42]<= -55; ws[7][2 ][43]<= -49; ws[7][2 ][44]<= -77; ws[7][2 ][45]<=-104; ws[7][2 ][46]<= -82; ws[7][2 ][47]<= -17; ws[7][2 ][48]<= -19;
        ws[7][3 ][0]<=  12; ws[7][3 ][1]<=  50; ws[7][3 ][2]<=  51; ws[7][3 ][3]<= 241; ws[7][3 ][4]<= 218; ws[7][3 ][5]<= 250; ws[7][3 ][6]<= 443; ws[7][3 ][7]<= -61; ws[7][3 ][8]<=  61; ws[7][3 ][9]<=  71; ws[7][3 ][10]<=  67; ws[7][3 ][11]<=  11; ws[7][3 ][12]<=  31; ws[7][3 ][13]<= 190; ws[7][3 ][14]<=   6; ws[7][3 ][15]<= 133; ws[7][3 ][16]<=  44; ws[7][3 ][17]<= -18; ws[7][3 ][18]<=  86; ws[7][3 ][19]<=  33; ws[7][3 ][20]<= 203; ws[7][3 ][21]<=  -6; ws[7][3 ][22]<=  98; ws[7][3 ][23]<=  29; ws[7][3 ][24]<=  28; ws[7][3 ][25]<= 172; ws[7][3 ][26]<=  45; ws[7][3 ][27]<= 278; ws[7][3 ][28]<=  -9; ws[7][3 ][29]<=  35; ws[7][3 ][30]<=  60; ws[7][3 ][31]<=  51; ws[7][3 ][32]<= 162; ws[7][3 ][33]<=   3; ws[7][3 ][34]<= 211; ws[7][3 ][35]<=   3; ws[7][3 ][36]<= -31; ws[7][3 ][37]<=  71; ws[7][3 ][38]<=   7; ws[7][3 ][39]<=  83; ws[7][3 ][40]<= -47; ws[7][3 ][41]<= 162; ws[7][3 ][42]<=  39; ws[7][3 ][43]<=  63; ws[7][3 ][44]<= 156; ws[7][3 ][45]<= 285; ws[7][3 ][46]<= 271; ws[7][3 ][47]<= 125; ws[7][3 ][48]<= 375;
        ws[7][4 ][0]<=  36; ws[7][4 ][1]<= 141; ws[7][4 ][2]<= 124; ws[7][4 ][3]<= -34; ws[7][4 ][4]<=  33; ws[7][4 ][5]<=  47; ws[7][4 ][6]<=  22; ws[7][4 ][7]<= -83; ws[7][4 ][8]<=  -4; ws[7][4 ][9]<= 214; ws[7][4 ][10]<=  47; ws[7][4 ][11]<=   2; ws[7][4 ][12]<=  33; ws[7][4 ][13]<=  -7; ws[7][4 ][14]<=-135; ws[7][4 ][15]<= -68; ws[7][4 ][16]<= 295; ws[7][4 ][17]<= -18; ws[7][4 ][18]<= -30; ws[7][4 ][19]<=  20; ws[7][4 ][20]<= -47; ws[7][4 ][21]<=-107; ws[7][4 ][22]<= -50; ws[7][4 ][23]<= 286; ws[7][4 ][24]<=   8; ws[7][4 ][25]<= -41; ws[7][4 ][26]<=  12; ws[7][4 ][27]<= -23; ws[7][4 ][28]<=-109; ws[7][4 ][29]<= -59; ws[7][4 ][30]<= 242; ws[7][4 ][31]<=   1; ws[7][4 ][32]<=   0; ws[7][4 ][33]<=  10; ws[7][4 ][34]<=  -5; ws[7][4 ][35]<= -96; ws[7][4 ][36]<= -29; ws[7][4 ][37]<= 134; ws[7][4 ][38]<= -52; ws[7][4 ][39]<=   1; ws[7][4 ][40]<=   9; ws[7][4 ][41]<= -21; ws[7][4 ][42]<=  24; ws[7][4 ][43]<= -30; ws[7][4 ][44]<=  40; ws[7][4 ][45]<=  12; ws[7][4 ][46]<=   2; ws[7][4 ][47]<= -11; ws[7][4 ][48]<= -82;
        ws[7][5 ][0]<=-172; ws[7][5 ][1]<=-156; ws[7][5 ][2]<=-106; ws[7][5 ][3]<=-158; ws[7][5 ][4]<=-187; ws[7][5 ][5]<= -69; ws[7][5 ][6]<=-207; ws[7][5 ][7]<=-145; ws[7][5 ][8]<=  10; ws[7][5 ][9]<=  15; ws[7][5 ][10]<=  12; ws[7][5 ][11]<=  15; ws[7][5 ][12]<=  42; ws[7][5 ][13]<= -58; ws[7][5 ][14]<=-130; ws[7][5 ][15]<= -13; ws[7][5 ][16]<=   7; ws[7][5 ][17]<= -15; ws[7][5 ][18]<= -31; ws[7][5 ][19]<=  38; ws[7][5 ][20]<= -24; ws[7][5 ][21]<= -85; ws[7][5 ][22]<=-112; ws[7][5 ][23]<= -55; ws[7][5 ][24]<= -70; ws[7][5 ][25]<= -65; ws[7][5 ][26]<= -17; ws[7][5 ][27]<= -10; ws[7][5 ][28]<= -82; ws[7][5 ][29]<= -81; ws[7][5 ][30]<= -21; ws[7][5 ][31]<=   0; ws[7][5 ][32]<= -50; ws[7][5 ][33]<=  21; ws[7][5 ][34]<= -17; ws[7][5 ][35]<= -23; ws[7][5 ][36]<= -39; ws[7][5 ][37]<= -40; ws[7][5 ][38]<=  32; ws[7][5 ][39]<= -16; ws[7][5 ][40]<=   5; ws[7][5 ][41]<=  -7; ws[7][5 ][42]<= -49; ws[7][5 ][43]<=-156; ws[7][5 ][44]<=-345; ws[7][5 ][45]<=-271; ws[7][5 ][46]<=-297; ws[7][5 ][47]<=-343; ws[7][5 ][48]<=-481;
        ws[7][6 ][0]<= 130; ws[7][6 ][1]<= -38; ws[7][6 ][2]<=  49; ws[7][6 ][3]<= 135; ws[7][6 ][4]<=  77; ws[7][6 ][5]<=   2; ws[7][6 ][6]<= -74; ws[7][6 ][7]<= -49; ws[7][6 ][8]<=-287; ws[7][6 ][9]<= -81; ws[7][6 ][10]<= -28; ws[7][6 ][11]<=   8; ws[7][6 ][12]<=  -8; ws[7][6 ][13]<= -97; ws[7][6 ][14]<= -79; ws[7][6 ][15]<=-219; ws[7][6 ][16]<=-212; ws[7][6 ][17]<= -72; ws[7][6 ][18]<= -12; ws[7][6 ][19]<= -58; ws[7][6 ][20]<= -75; ws[7][6 ][21]<=  12; ws[7][6 ][22]<=-124; ws[7][6 ][23]<=-188; ws[7][6 ][24]<=-118; ws[7][6 ][25]<=   4; ws[7][6 ][26]<= -87; ws[7][6 ][27]<= -80; ws[7][6 ][28]<=  -4; ws[7][6 ][29]<= -69; ws[7][6 ][30]<=-106; ws[7][6 ][31]<= -83; ws[7][6 ][32]<= -14; ws[7][6 ][33]<= -96; ws[7][6 ][34]<= -52; ws[7][6 ][35]<=  19; ws[7][6 ][36]<=  20; ws[7][6 ][37]<= -17; ws[7][6 ][38]<=  70; ws[7][6 ][39]<=  -8; ws[7][6 ][40]<= -51; ws[7][6 ][41]<=   2; ws[7][6 ][42]<=  26; ws[7][6 ][43]<=  28; ws[7][6 ][44]<= -73; ws[7][6 ][45]<= -36; ws[7][6 ][46]<= 104; ws[7][6 ][47]<= -52; ws[7][6 ][48]<=  -6;
        ws[7][7 ][0]<=-101; ws[7][7 ][1]<= -31; ws[7][7 ][2]<= -57; ws[7][7 ][3]<= -22; ws[7][7 ][4]<= 107; ws[7][7 ][5]<= 147; ws[7][7 ][6]<= 178; ws[7][7 ][7]<= -76; ws[7][7 ][8]<= -42; ws[7][7 ][9]<= -65; ws[7][7 ][10]<= -44; ws[7][7 ][11]<=  36; ws[7][7 ][12]<= 101; ws[7][7 ][13]<= 166; ws[7][7 ][14]<= -11; ws[7][7 ][15]<= -40; ws[7][7 ][16]<= -70; ws[7][7 ][17]<= -37; ws[7][7 ][18]<=  -9; ws[7][7 ][19]<=  39; ws[7][7 ][20]<= 137; ws[7][7 ][21]<=  -4; ws[7][7 ][22]<= -14; ws[7][7 ][23]<=  -2; ws[7][7 ][24]<= -49; ws[7][7 ][25]<=   6; ws[7][7 ][26]<= -30; ws[7][7 ][27]<= 144; ws[7][7 ][28]<=  -7; ws[7][7 ][29]<=  79; ws[7][7 ][30]<=  90; ws[7][7 ][31]<= -37; ws[7][7 ][32]<= -76; ws[7][7 ][33]<=  18; ws[7][7 ][34]<= 111; ws[7][7 ][35]<=  65; ws[7][7 ][36]<=  86; ws[7][7 ][37]<=  80; ws[7][7 ][38]<=-126; ws[7][7 ][39]<= -61; ws[7][7 ][40]<= -15; ws[7][7 ][41]<= 115; ws[7][7 ][42]<=  44; ws[7][7 ][43]<= -26; ws[7][7 ][44]<=   5; ws[7][7 ][45]<= -18; ws[7][7 ][46]<= -12; ws[7][7 ][47]<=  59; ws[7][7 ][48]<= 106;
        ws[7][8 ][0]<= -62; ws[7][8 ][1]<=-132; ws[7][8 ][2]<=-228; ws[7][8 ][3]<=-108; ws[7][8 ][4]<=-134; ws[7][8 ][5]<=-326; ws[7][8 ][6]<=-285; ws[7][8 ][7]<=   9; ws[7][8 ][8]<= -62; ws[7][8 ][9]<=-145; ws[7][8 ][10]<=  34; ws[7][8 ][11]<=  26; ws[7][8 ][12]<=  -3; ws[7][8 ][13]<=-104; ws[7][8 ][14]<= -77; ws[7][8 ][15]<= -95; ws[7][8 ][16]<= -43; ws[7][8 ][17]<=-133; ws[7][8 ][18]<=  30; ws[7][8 ][19]<=  50; ws[7][8 ][20]<=-102; ws[7][8 ][21]<= -18; ws[7][8 ][22]<= -51; ws[7][8 ][23]<=-190; ws[7][8 ][24]<=-227; ws[7][8 ][25]<=  91; ws[7][8 ][26]<= -31; ws[7][8 ][27]<= -57; ws[7][8 ][28]<=  45; ws[7][8 ][29]<=  66; ws[7][8 ][30]<=-151; ws[7][8 ][31]<=-192; ws[7][8 ][32]<= 167; ws[7][8 ][33]<= -44; ws[7][8 ][34]<=  84; ws[7][8 ][35]<=  37; ws[7][8 ][36]<=  35; ws[7][8 ][37]<= -32; ws[7][8 ][38]<= -58; ws[7][8 ][39]<= 156; ws[7][8 ][40]<= -88; ws[7][8 ][41]<=  81; ws[7][8 ][42]<= -17; ws[7][8 ][43]<= -28; ws[7][8 ][44]<= -15; ws[7][8 ][45]<=-213; ws[7][8 ][46]<=  59; ws[7][8 ][47]<= -32; ws[7][8 ][48]<= -26;
        ws[7][9 ][0]<=  61; ws[7][9 ][1]<=  -7; ws[7][9 ][2]<= 136; ws[7][9 ][3]<= 205; ws[7][9 ][4]<= 184; ws[7][9 ][5]<=  51; ws[7][9 ][6]<= -13; ws[7][9 ][7]<=   3; ws[7][9 ][8]<=  66; ws[7][9 ][9]<= 163; ws[7][9 ][10]<= 173; ws[7][9 ][11]<= 117; ws[7][9 ][12]<= -31; ws[7][9 ][13]<=   3; ws[7][9 ][14]<=  37; ws[7][9 ][15]<=  96; ws[7][9 ][16]<=  69; ws[7][9 ][17]<=  72; ws[7][9 ][18]<= 108; ws[7][9 ][19]<=  -4; ws[7][9 ][20]<=  21; ws[7][9 ][21]<=  37; ws[7][9 ][22]<=  59; ws[7][9 ][23]<=   6; ws[7][9 ][24]<= 105; ws[7][9 ][25]<=  62; ws[7][9 ][26]<= -16; ws[7][9 ][27]<=  20; ws[7][9 ][28]<= -45; ws[7][9 ][29]<=  -5; ws[7][9 ][30]<=  63; ws[7][9 ][31]<=  39; ws[7][9 ][32]<=  69; ws[7][9 ][33]<=  12; ws[7][9 ][34]<=  -8; ws[7][9 ][35]<=  -9; ws[7][9 ][36]<=  12; ws[7][9 ][37]<= 175; ws[7][9 ][38]<=  83; ws[7][9 ][39]<=  28; ws[7][9 ][40]<= -28; ws[7][9 ][41]<=  17; ws[7][9 ][42]<=  14; ws[7][9 ][43]<=  13; ws[7][9 ][44]<= 169; ws[7][9 ][45]<= 110; ws[7][9 ][46]<=  60; ws[7][9 ][47]<= -17; ws[7][9 ][48]<=   3;
        ws[7][10][0]<= -93; ws[7][10][1]<= -83; ws[7][10][2]<=   5; ws[7][10][3]<= -90; ws[7][10][4]<=-166; ws[7][10][5]<=-145; ws[7][10][6]<=-163; ws[7][10][7]<=  21; ws[7][10][8]<=-114; ws[7][10][9]<=  -5; ws[7][10][10]<=-120; ws[7][10][11]<= -95; ws[7][10][12]<= -77; ws[7][10][13]<=-183; ws[7][10][14]<=  28; ws[7][10][15]<= -84; ws[7][10][16]<=  33; ws[7][10][17]<= -82; ws[7][10][18]<= -28; ws[7][10][19]<= -17; ws[7][10][20]<= -89; ws[7][10][21]<=  40; ws[7][10][22]<= -97; ws[7][10][23]<= -21; ws[7][10][24]<= -19; ws[7][10][25]<= -61; ws[7][10][26]<=  30; ws[7][10][27]<=-119; ws[7][10][28]<= -53; ws[7][10][29]<= -90; ws[7][10][30]<=   3; ws[7][10][31]<= -68; ws[7][10][32]<= -71; ws[7][10][33]<= -77; ws[7][10][34]<=-122; ws[7][10][35]<= -66; ws[7][10][36]<=-115; ws[7][10][37]<= -73; ws[7][10][38]<= -65; ws[7][10][39]<= -89; ws[7][10][40]<=-125; ws[7][10][41]<=-113; ws[7][10][42]<=  -3; ws[7][10][43]<=-104; ws[7][10][44]<= -88; ws[7][10][45]<=-105; ws[7][10][46]<= -67; ws[7][10][47]<=-123; ws[7][10][48]<=-197;
        ws[7][11][0]<= -55; ws[7][11][1]<=  34; ws[7][11][2]<= 107; ws[7][11][3]<= 123; ws[7][11][4]<= 148; ws[7][11][5]<= 100; ws[7][11][6]<= 166; ws[7][11][7]<= -37; ws[7][11][8]<=  59; ws[7][11][9]<= 112; ws[7][11][10]<= 121; ws[7][11][11]<= 131; ws[7][11][12]<= 127; ws[7][11][13]<= 120; ws[7][11][14]<=  32; ws[7][11][15]<=  64; ws[7][11][16]<=  92; ws[7][11][17]<=  83; ws[7][11][18]<=  63; ws[7][11][19]<= 114; ws[7][11][20]<=  70; ws[7][11][21]<=  26; ws[7][11][22]<=  57; ws[7][11][23]<= 118; ws[7][11][24]<= 127; ws[7][11][25]<= 114; ws[7][11][26]<=  83; ws[7][11][27]<=  18; ws[7][11][28]<=  73; ws[7][11][29]<=  81; ws[7][11][30]<= 161; ws[7][11][31]<=  89; ws[7][11][32]<=  50; ws[7][11][33]<=  85; ws[7][11][34]<= -40; ws[7][11][35]<=  90; ws[7][11][36]<= 134; ws[7][11][37]<= 155; ws[7][11][38]<=  71; ws[7][11][39]<=  56; ws[7][11][40]<=  78; ws[7][11][41]<= -46; ws[7][11][42]<= 110; ws[7][11][43]<= 109; ws[7][11][44]<= 165; ws[7][11][45]<=  87; ws[7][11][46]<= 134; ws[7][11][47]<=  97; ws[7][11][48]<=   3;
        ws[7][12][0]<= -23; ws[7][12][1]<=  22; ws[7][12][2]<=  18; ws[7][12][3]<= 115; ws[7][12][4]<= 122; ws[7][12][5]<=  51; ws[7][12][6]<=  67; ws[7][12][7]<= -31; ws[7][12][8]<= -23; ws[7][12][9]<= -25; ws[7][12][10]<=  20; ws[7][12][11]<= 100; ws[7][12][12]<= -26; ws[7][12][13]<=  19; ws[7][12][14]<= -67; ws[7][12][15]<=   0; ws[7][12][16]<= -77; ws[7][12][17]<= -36; ws[7][12][18]<= 139; ws[7][12][19]<=  74; ws[7][12][20]<=  29; ws[7][12][21]<=  61; ws[7][12][22]<=  -5; ws[7][12][23]<= -16; ws[7][12][24]<=-113; ws[7][12][25]<=  56; ws[7][12][26]<=  51; ws[7][12][27]<=  41; ws[7][12][28]<=  51; ws[7][12][29]<= -25; ws[7][12][30]<= -24; ws[7][12][31]<=-128; ws[7][12][32]<=  19; ws[7][12][33]<=  89; ws[7][12][34]<=  82; ws[7][12][35]<=  48; ws[7][12][36]<= -53; ws[7][12][37]<=  -6; ws[7][12][38]<= -75; ws[7][12][39]<=  23; ws[7][12][40]<= 166; ws[7][12][41]<= 112; ws[7][12][42]<=  93; ws[7][12][43]<=  80; ws[7][12][44]<= 153; ws[7][12][45]<=  46; ws[7][12][46]<=   1; ws[7][12][47]<=  93; ws[7][12][48]<= 182;
        ws[7][13][0]<= -43; ws[7][13][1]<=-227; ws[7][13][2]<=-234; ws[7][13][3]<=-187; ws[7][13][4]<=  26; ws[7][13][5]<=  -2; ws[7][13][6]<=-219; ws[7][13][7]<= -38; ws[7][13][8]<= -37; ws[7][13][9]<=-191; ws[7][13][10]<= -48; ws[7][13][11]<=  94; ws[7][13][12]<= -11; ws[7][13][13]<=-108; ws[7][13][14]<=   8; ws[7][13][15]<=  14; ws[7][13][16]<=-206; ws[7][13][17]<=  29; ws[7][13][18]<=  36; ws[7][13][19]<=  34; ws[7][13][20]<= -16; ws[7][13][21]<=  42; ws[7][13][22]<=  13; ws[7][13][23]<=-141; ws[7][13][24]<=  12; ws[7][13][25]<=  48; ws[7][13][26]<= 112; ws[7][13][27]<= 113; ws[7][13][28]<=  45; ws[7][13][29]<= -55; ws[7][13][30]<=-163; ws[7][13][31]<=   4; ws[7][13][32]<=  46; ws[7][13][33]<=  98; ws[7][13][34]<= 132; ws[7][13][35]<= -26; ws[7][13][36]<= -83; ws[7][13][37]<= -79; ws[7][13][38]<=  56; ws[7][13][39]<=  32; ws[7][13][40]<=  85; ws[7][13][41]<=  68; ws[7][13][42]<= -62; ws[7][13][43]<=-147; ws[7][13][44]<= -72; ws[7][13][45]<=  38; ws[7][13][46]<= -29; ws[7][13][47]<= -86; ws[7][13][48]<=  43;
        ws[7][14][0]<= -10; ws[7][14][1]<= 210; ws[7][14][2]<=  -3; ws[7][14][3]<=-148; ws[7][14][4]<=-230; ws[7][14][5]<= -39; ws[7][14][6]<= -68; ws[7][14][7]<= -68; ws[7][14][8]<= 137; ws[7][14][9]<= -30; ws[7][14][10]<=-109; ws[7][14][11]<= -84; ws[7][14][12]<= -30; ws[7][14][13]<= -19; ws[7][14][14]<=-128; ws[7][14][15]<=  15; ws[7][14][16]<= -34; ws[7][14][17]<= -38; ws[7][14][18]<= -40; ws[7][14][19]<=  32; ws[7][14][20]<=  19; ws[7][14][21]<=-253; ws[7][14][22]<= -47; ws[7][14][23]<=   3; ws[7][14][24]<=   9; ws[7][14][25]<= -20; ws[7][14][26]<= -45; ws[7][14][27]<=  17; ws[7][14][28]<=-213; ws[7][14][29]<= -64; ws[7][14][30]<=  -9; ws[7][14][31]<=   4; ws[7][14][32]<= -59; ws[7][14][33]<= -90; ws[7][14][34]<= -66; ws[7][14][35]<=-146; ws[7][14][36]<=  -4; ws[7][14][37]<= -62; ws[7][14][38]<=-128; ws[7][14][39]<= -59; ws[7][14][40]<=-192; ws[7][14][41]<= -61; ws[7][14][42]<= -42; ws[7][14][43]<=-141; ws[7][14][44]<=-121; ws[7][14][45]<=-105; ws[7][14][46]<=-130; ws[7][14][47]<=-249; ws[7][14][48]<=-251;
        ws[7][15][0]<=-262; ws[7][15][1]<=-256; ws[7][15][2]<=-224; ws[7][15][3]<= -83; ws[7][15][4]<=  18; ws[7][15][5]<=  27; ws[7][15][6]<= -69; ws[7][15][7]<=-127; ws[7][15][8]<=-147; ws[7][15][9]<= -69; ws[7][15][10]<= -26; ws[7][15][11]<=  38; ws[7][15][12]<=  56; ws[7][15][13]<=  13; ws[7][15][14]<= -65; ws[7][15][15]<=-107; ws[7][15][16]<= -40; ws[7][15][17]<= -80; ws[7][15][18]<=  -3; ws[7][15][19]<=   2; ws[7][15][20]<= -71; ws[7][15][21]<= -91; ws[7][15][22]<=  24; ws[7][15][23]<=  39; ws[7][15][24]<= -39; ws[7][15][25]<= -43; ws[7][15][26]<= -54; ws[7][15][27]<=   2; ws[7][15][28]<= -90; ws[7][15][29]<= -31; ws[7][15][30]<=-120; ws[7][15][31]<=-141; ws[7][15][32]<=-110; ws[7][15][33]<= -19; ws[7][15][34]<=   1; ws[7][15][35]<=-113; ws[7][15][36]<=-120; ws[7][15][37]<=-215; ws[7][15][38]<=-136; ws[7][15][39]<= -80; ws[7][15][40]<=  24; ws[7][15][41]<=  24; ws[7][15][42]<=-261; ws[7][15][43]<=-137; ws[7][15][44]<=-120; ws[7][15][45]<= -60; ws[7][15][46]<=-130; ws[7][15][47]<= -83; ws[7][15][48]<= -54;
    end

    always@(posedge clk) begin
        if(rst) begin
            w0 <=0; w1 <=0; w2 <=0; w3 <=0; w4 <=0; w5 <=0; w6 <=0;
            w7 <=0; w8 <=0; w9 <=0; w10<=0; w11<=0; w12<=0; w13<=0;
            w14<=0; w15<=0; w16<=0; w17<=0; w18<=0; w19<=0; w20<=0;
            w21<=0; w22<=0; w23<=0; w24<=0; w25<=0; w26<=0; w27<=0;
            w28<=0; w29<=0; w30<=0; w31<=0; w32<=0; w33<=0; w34<=0;
            w35<=0; w36<=0; w37<=0; w38<=0; w39<=0; w40<=0; w41<=0;
            w42<=0; w43<=0; w44<=0; w45<=0; w46<=0; w47<=0; w48<=0;
            ready<=0;
        end else if(start) begin
            w0 <=ws[layer_sel][filter_sel][0 ]; w1 <=ws[layer_sel][filter_sel][1 ]; w2 <=ws[layer_sel][filter_sel][2 ]; w3 <=ws[layer_sel][filter_sel][3 ]; w4 <=ws[layer_sel][filter_sel][4 ]; w5 <=ws[layer_sel][filter_sel][5 ]; w6 <=ws[layer_sel][filter_sel][6 ];
            w7 <=ws[layer_sel][filter_sel][7 ]; w8 <=ws[layer_sel][filter_sel][8 ]; w9 <=ws[layer_sel][filter_sel][9 ]; w10<=ws[layer_sel][filter_sel][10]; w11<=ws[layer_sel][filter_sel][11]; w12<=ws[layer_sel][filter_sel][12]; w13<=ws[layer_sel][filter_sel][13];
            w14<=ws[layer_sel][filter_sel][14]; w15<=ws[layer_sel][filter_sel][15]; w16<=ws[layer_sel][filter_sel][16]; w17<=ws[layer_sel][filter_sel][17]; w18<=ws[layer_sel][filter_sel][18]; w19<=ws[layer_sel][filter_sel][19]; w20<=ws[layer_sel][filter_sel][20];
            w21<=ws[layer_sel][filter_sel][21]; w22<=ws[layer_sel][filter_sel][22]; w23<=ws[layer_sel][filter_sel][23]; w24<=ws[layer_sel][filter_sel][24]; w25<=ws[layer_sel][filter_sel][25]; w26<=ws[layer_sel][filter_sel][26]; w27<=ws[layer_sel][filter_sel][27];
            w28<=ws[layer_sel][filter_sel][28]; w29<=ws[layer_sel][filter_sel][29]; w30<=ws[layer_sel][filter_sel][30]; w31<=ws[layer_sel][filter_sel][31]; w32<=ws[layer_sel][filter_sel][32]; w33<=ws[layer_sel][filter_sel][33]; w34<=ws[layer_sel][filter_sel][34];
            w35<=ws[layer_sel][filter_sel][35]; w36<=ws[layer_sel][filter_sel][36]; w37<=ws[layer_sel][filter_sel][37]; w38<=ws[layer_sel][filter_sel][38]; w39<=ws[layer_sel][filter_sel][39]; w40<=ws[layer_sel][filter_sel][40]; w41<=ws[layer_sel][filter_sel][41];
            w42<=ws[layer_sel][filter_sel][42]; w43<=ws[layer_sel][filter_sel][43]; w44<=ws[layer_sel][filter_sel][44]; w45<=ws[layer_sel][filter_sel][45]; w46<=ws[layer_sel][filter_sel][46]; w47<=ws[layer_sel][filter_sel][47]; w48<=ws[layer_sel][filter_sel][48];
            ready<=1;
        end
    end
endmodule