`timescale 1ns/ 1ps

module dsconv_block_pointwise_weights_memory(
    input  wire                clk,
    input  wire                rst,
    input  wire                start,
    input  wire        [2: 0]  layer_sel,     // 8
    input  wire        [3: 0]  input_filter,  // 16
    input  wire        [3: 0]  output_filter, // 16
    output reg  signed [17: 0] w,
    output reg                 ready
);
    reg signed [17: 0] ws [0: 7][0: 15][0: 15];

    initial begin
        ws[0][0 ][0]<=  83; ws[0][0 ][1]<=-438; ws[0][0 ][2]<=  49; ws[0][0 ][3]<=  97; ws[0][0 ][4]<=-149; ws[0][0 ][5]<= 150; ws[0][0 ][6]<=  68; ws[0][0 ][7]<=-217; ws[0][0 ][8]<= 155; ws[0][0 ][9]<=-133; ws[0][0 ][10]<=-331; ws[0][0 ][11]<= 138; ws[0][0 ][12]<= 199; ws[0][0 ][13]<= -24; ws[0][0 ][14]<=  92; ws[0][0 ][15]<=-130;
        ws[0][1 ][0]<=  56; ws[0][1 ][1]<=  72; ws[0][1 ][2]<=  30; ws[0][1 ][3]<= 125; ws[0][1 ][4]<=-219; ws[0][1 ][5]<= 182; ws[0][1 ][6]<=  38; ws[0][1 ][7]<= -66; ws[0][1 ][8]<= 280; ws[0][1 ][9]<=-147; ws[0][1 ][10]<= 366; ws[0][1 ][11]<= -72; ws[0][1 ][12]<=-251; ws[0][1 ][13]<= -55; ws[0][1 ][14]<=  34; ws[0][1 ][15]<=  48;
        ws[0][2 ][0]<= 299; ws[0][2 ][1]<=  81; ws[0][2 ][2]<=  98; ws[0][2 ][3]<= 235; ws[0][2 ][4]<=  -9; ws[0][2 ][5]<= -11; ws[0][2 ][6]<= 213; ws[0][2 ][7]<= 244; ws[0][2 ][8]<= 150; ws[0][2 ][9]<=  56; ws[0][2 ][10]<= 128; ws[0][2 ][11]<=-113; ws[0][2 ][12]<=  42; ws[0][2 ][13]<=   3; ws[0][2 ][14]<=  67; ws[0][2 ][15]<= 432;
        ws[0][3 ][0]<= -65; ws[0][3 ][1]<= 184; ws[0][3 ][2]<=-102; ws[0][3 ][3]<= 420; ws[0][3 ][4]<=-236; ws[0][3 ][5]<=  -5; ws[0][3 ][6]<=   9; ws[0][3 ][7]<=  90; ws[0][3 ][8]<=-353; ws[0][3 ][9]<=  32; ws[0][3 ][10]<= 223; ws[0][3 ][11]<= -58; ws[0][3 ][12]<= -54; ws[0][3 ][13]<= 332; ws[0][3 ][14]<=  53; ws[0][3 ][15]<=  27;
        ws[0][4 ][0]<= -42; ws[0][4 ][1]<=-194; ws[0][4 ][2]<=-147; ws[0][4 ][3]<= 107; ws[0][4 ][4]<= 123; ws[0][4 ][5]<= 192; ws[0][4 ][6]<= -61; ws[0][4 ][7]<=-123; ws[0][4 ][8]<= 169; ws[0][4 ][9]<= 386; ws[0][4 ][10]<=-135; ws[0][4 ][11]<= 157; ws[0][4 ][12]<= 397; ws[0][4 ][13]<=-189; ws[0][4 ][14]<=   7; ws[0][4 ][15]<=  40;
        ws[0][5 ][0]<=  44; ws[0][5 ][1]<=-151; ws[0][5 ][2]<= 144; ws[0][5 ][3]<=-254; ws[0][5 ][4]<=-107; ws[0][5 ][5]<=-247; ws[0][5 ][6]<= 115; ws[0][5 ][7]<=-278; ws[0][5 ][8]<=  18; ws[0][5 ][9]<= -93; ws[0][5 ][10]<=  70; ws[0][5 ][11]<=-233; ws[0][5 ][12]<= -98; ws[0][5 ][13]<=   6; ws[0][5 ][14]<=-324; ws[0][5 ][15]<=  13;
        ws[0][6 ][0]<=-250; ws[0][6 ][1]<=  33; ws[0][6 ][2]<=   9; ws[0][6 ][3]<=-204; ws[0][6 ][4]<= -10; ws[0][6 ][5]<=  19; ws[0][6 ][6]<=-793; ws[0][6 ][7]<=-195; ws[0][6 ][8]<= -40; ws[0][6 ][9]<= -71; ws[0][6 ][10]<=  44; ws[0][6 ][11]<= 230; ws[0][6 ][12]<= -55; ws[0][6 ][13]<=  81; ws[0][6 ][14]<=-182; ws[0][6 ][15]<=  -7;
        ws[0][7 ][0]<= 121; ws[0][7 ][1]<=-110; ws[0][7 ][2]<=-325; ws[0][7 ][3]<=  23; ws[0][7 ][4]<=-264; ws[0][7 ][5]<=-204; ws[0][7 ][6]<= -23; ws[0][7 ][7]<= 108; ws[0][7 ][8]<= 284; ws[0][7 ][9]<= 257; ws[0][7 ][10]<=-151; ws[0][7 ][11]<=  14; ws[0][7 ][12]<= 213; ws[0][7 ][13]<= -53; ws[0][7 ][14]<=-235; ws[0][7 ][15]<= -72;
        ws[0][8 ][0]<= 343; ws[0][8 ][1]<=  32; ws[0][8 ][2]<=-218; ws[0][8 ][3]<=-105; ws[0][8 ][4]<=  85; ws[0][8 ][5]<=-139; ws[0][8 ][6]<=  45; ws[0][8 ][7]<=-121; ws[0][8 ][8]<=-163; ws[0][8 ][9]<=  39; ws[0][8 ][10]<= -14; ws[0][8 ][11]<=  68; ws[0][8 ][12]<= 261; ws[0][8 ][13]<=  -5; ws[0][8 ][14]<= -50; ws[0][8 ][15]<= 184;
        ws[0][9 ][0]<= 197; ws[0][9 ][1]<=  81; ws[0][9 ][2]<=  18; ws[0][9 ][3]<= 124; ws[0][9 ][4]<= 124; ws[0][9 ][5]<=-133; ws[0][9 ][6]<=-150; ws[0][9 ][7]<=  -1; ws[0][9 ][8]<=-182; ws[0][9 ][9]<= -63; ws[0][9 ][10]<= -62; ws[0][9 ][11]<=-172; ws[0][9 ][12]<=  40; ws[0][9 ][13]<=-422; ws[0][9 ][14]<= -39; ws[0][9 ][15]<=-353;
        ws[0][10][0]<=  95; ws[0][10][1]<=-214; ws[0][10][2]<=  51; ws[0][10][3]<= 205; ws[0][10][4]<=   7; ws[0][10][5]<=-223; ws[0][10][6]<= -78; ws[0][10][7]<=  39; ws[0][10][8]<=-105; ws[0][10][9]<= -90; ws[0][10][10]<= 183; ws[0][10][11]<=-124; ws[0][10][12]<= 158; ws[0][10][13]<= 188; ws[0][10][14]<= -53; ws[0][10][15]<= -76;
        ws[0][11][0]<=  -1; ws[0][11][1]<= 121; ws[0][11][2]<= 147; ws[0][11][3]<=-216; ws[0][11][4]<=-183; ws[0][11][5]<=-105; ws[0][11][6]<= -69; ws[0][11][7]<=  87; ws[0][11][8]<= 197; ws[0][11][9]<= 156; ws[0][11][10]<= 364; ws[0][11][11]<=  17; ws[0][11][12]<=-160; ws[0][11][13]<= 212; ws[0][11][14]<= -80; ws[0][11][15]<= -39;
        ws[0][12][0]<=-100; ws[0][12][1]<=-351; ws[0][12][2]<=-175; ws[0][12][3]<= 377; ws[0][12][4]<=  54; ws[0][12][5]<= 506; ws[0][12][6]<= -82; ws[0][12][7]<= 189; ws[0][12][8]<=  61; ws[0][12][9]<=-176; ws[0][12][10]<= 124; ws[0][12][11]<=-378; ws[0][12][12]<=-176; ws[0][12][13]<= 422; ws[0][12][14]<= 303; ws[0][12][15]<= 139;
        ws[0][13][0]<= -37; ws[0][13][1]<= 162; ws[0][13][2]<=  62; ws[0][13][3]<=-257; ws[0][13][4]<=  78; ws[0][13][5]<= 174; ws[0][13][6]<=  60; ws[0][13][7]<=-192; ws[0][13][8]<= 206; ws[0][13][9]<= -92; ws[0][13][10]<=  30; ws[0][13][11]<= -25; ws[0][13][12]<= 120; ws[0][13][13]<=-218; ws[0][13][14]<=  14; ws[0][13][15]<=  31;
        ws[0][14][0]<= -18; ws[0][14][1]<=  49; ws[0][14][2]<= 184; ws[0][14][3]<=-117; ws[0][14][4]<=-400; ws[0][14][5]<=-129; ws[0][14][6]<= 103; ws[0][14][7]<=-213; ws[0][14][8]<=-182; ws[0][14][9]<= 126; ws[0][14][10]<= 158; ws[0][14][11]<=  28; ws[0][14][12]<= 122; ws[0][14][13]<=  37; ws[0][14][14]<= -41; ws[0][14][15]<=-112;
        ws[0][15][0]<= 157; ws[0][15][1]<= 209; ws[0][15][2]<=  31; ws[0][15][3]<= -78; ws[0][15][4]<= -91; ws[0][15][5]<= 197; ws[0][15][6]<= 106; ws[0][15][7]<=-271; ws[0][15][8]<=-213; ws[0][15][9]<=  96; ws[0][15][10]<=  83; ws[0][15][11]<=-162; ws[0][15][12]<= 108; ws[0][15][13]<=  39; ws[0][15][14]<= -51; ws[0][15][15]<= -61;

        ws[1][0 ][0]<=-211; ws[1][0 ][1]<= -59; ws[1][0 ][2]<= 182; ws[1][0 ][3]<= -43; ws[1][0 ][4]<= 177; ws[1][0 ][5]<= -79; ws[1][0 ][6]<=-171; ws[1][0 ][7]<= -87; ws[1][0 ][8]<=  89; ws[1][0 ][9]<= 262; ws[1][0 ][10]<= -15; ws[1][0 ][11]<= -52; ws[1][0 ][12]<= -65; ws[1][0 ][13]<= 164; ws[1][0 ][14]<=  71; ws[1][0 ][15]<= -11;
        ws[1][1 ][0]<=  62; ws[1][1 ][1]<=  42; ws[1][1 ][2]<= -15; ws[1][1 ][3]<= -71; ws[1][1 ][4]<= -20; ws[1][1 ][5]<=  50; ws[1][1 ][6]<= -37; ws[1][1 ][7]<=   2; ws[1][1 ][8]<=  77; ws[1][1 ][9]<= 111; ws[1][1 ][10]<=  23; ws[1][1 ][11]<= -75; ws[1][1 ][12]<=-461; ws[1][1 ][13]<=  65; ws[1][1 ][14]<=-154; ws[1][1 ][15]<= 395;
        ws[1][2 ][0]<=-340; ws[1][2 ][1]<=-139; ws[1][2 ][2]<=-170; ws[1][2 ][3]<=-152; ws[1][2 ][4]<= -62; ws[1][2 ][5]<=-351; ws[1][2 ][6]<= 187; ws[1][2 ][7]<=-145; ws[1][2 ][8]<= 110; ws[1][2 ][9]<=-107; ws[1][2 ][10]<= 104; ws[1][2 ][11]<=-115; ws[1][2 ][12]<= 261; ws[1][2 ][13]<= 227; ws[1][2 ][14]<= -24; ws[1][2 ][15]<=   2;
        ws[1][3 ][0]<=  37; ws[1][3 ][1]<= 152; ws[1][3 ][2]<= 209; ws[1][3 ][3]<=  80; ws[1][3 ][4]<= 156; ws[1][3 ][5]<=-117; ws[1][3 ][6]<=  48; ws[1][3 ][7]<= 148; ws[1][3 ][8]<=  15; ws[1][3 ][9]<= -29; ws[1][3 ][10]<= 110; ws[1][3 ][11]<=  71; ws[1][3 ][12]<=-192; ws[1][3 ][13]<= 229; ws[1][3 ][14]<=-190; ws[1][3 ][15]<=-100;
        ws[1][4 ][0]<= -80; ws[1][4 ][1]<=  69; ws[1][4 ][2]<= 289; ws[1][4 ][3]<= 126; ws[1][4 ][4]<=  43; ws[1][4 ][5]<=  24; ws[1][4 ][6]<= 162; ws[1][4 ][7]<=-124; ws[1][4 ][8]<= 357; ws[1][4 ][9]<= -98; ws[1][4 ][10]<= 174; ws[1][4 ][11]<=-126; ws[1][4 ][12]<=-132; ws[1][4 ][13]<=-116; ws[1][4 ][14]<=-296; ws[1][4 ][15]<= -37;
        ws[1][5 ][0]<=-234; ws[1][5 ][1]<= 112; ws[1][5 ][2]<= 131; ws[1][5 ][3]<=  46; ws[1][5 ][4]<=  72; ws[1][5 ][5]<= -52; ws[1][5 ][6]<=-225; ws[1][5 ][7]<=-313; ws[1][5 ][8]<=-110; ws[1][5 ][9]<=-104; ws[1][5 ][10]<=-173; ws[1][5 ][11]<=-369; ws[1][5 ][12]<=-113; ws[1][5 ][13]<=  36; ws[1][5 ][14]<= 296; ws[1][5 ][15]<= -86;
        ws[1][6 ][0]<=  59; ws[1][6 ][1]<=  54; ws[1][6 ][2]<= -18; ws[1][6 ][3]<=-149; ws[1][6 ][4]<= 517; ws[1][6 ][5]<= -34; ws[1][6 ][6]<= 133; ws[1][6 ][7]<= -46; ws[1][6 ][8]<=  -6; ws[1][6 ][9]<= 285; ws[1][6 ][10]<= 267; ws[1][6 ][11]<=   4; ws[1][6 ][12]<=  26; ws[1][6 ][13]<= -48; ws[1][6 ][14]<= -84; ws[1][6 ][15]<= -48;
        ws[1][7 ][0]<=-165; ws[1][7 ][1]<= -59; ws[1][7 ][2]<=-115; ws[1][7 ][3]<= -71; ws[1][7 ][4]<= 256; ws[1][7 ][5]<=  32; ws[1][7 ][6]<=   6; ws[1][7 ][7]<= 158; ws[1][7 ][8]<=-242; ws[1][7 ][9]<=-222; ws[1][7 ][10]<=  32; ws[1][7 ][11]<= -51; ws[1][7 ][12]<= -39; ws[1][7 ][13]<= 105; ws[1][7 ][14]<=-157; ws[1][7 ][15]<=-133;
        ws[1][8 ][0]<= 314; ws[1][8 ][1]<= 345; ws[1][8 ][2]<=-126; ws[1][8 ][3]<= 167; ws[1][8 ][4]<=  -2; ws[1][8 ][5]<= 303; ws[1][8 ][6]<=-194; ws[1][8 ][7]<=   5; ws[1][8 ][8]<=-163; ws[1][8 ][9]<=  61; ws[1][8 ][10]<= 222; ws[1][8 ][11]<=  27; ws[1][8 ][12]<= 146; ws[1][8 ][13]<=-110; ws[1][8 ][14]<= -79; ws[1][8 ][15]<= 215;
        ws[1][9 ][0]<=  30; ws[1][9 ][1]<=  -7; ws[1][9 ][2]<= -71; ws[1][9 ][3]<= 411; ws[1][9 ][4]<= -33; ws[1][9 ][5]<= 269; ws[1][9 ][6]<=  25; ws[1][9 ][7]<= 236; ws[1][9 ][8]<=-337; ws[1][9 ][9]<= 103; ws[1][9 ][10]<=  47; ws[1][9 ][11]<= -81; ws[1][9 ][12]<= 223; ws[1][9 ][13]<= 183; ws[1][9 ][14]<=-293; ws[1][9 ][15]<=-315;
        ws[1][10][0]<= 192; ws[1][10][1]<= 103; ws[1][10][2]<=-173; ws[1][10][3]<=-125; ws[1][10][4]<=  45; ws[1][10][5]<= 309; ws[1][10][6]<=-237; ws[1][10][7]<= -40; ws[1][10][8]<=  51; ws[1][10][9]<= 204; ws[1][10][10]<= 143; ws[1][10][11]<= 184; ws[1][10][12]<= -24; ws[1][10][13]<= -63; ws[1][10][14]<= -88; ws[1][10][15]<=  55;
        ws[1][11][0]<=-242; ws[1][11][1]<=-274; ws[1][11][2]<= 249; ws[1][11][3]<= 112; ws[1][11][4]<= -85; ws[1][11][5]<=-207; ws[1][11][6]<= 171; ws[1][11][7]<= 241; ws[1][11][8]<= -52; ws[1][11][9]<= -39; ws[1][11][10]<= -99; ws[1][11][11]<= 117; ws[1][11][12]<= -10; ws[1][11][13]<= 232; ws[1][11][14]<= 173; ws[1][11][15]<=  78;
        ws[1][12][0]<=  -7; ws[1][12][1]<=  12; ws[1][12][2]<= 220; ws[1][12][3]<= -40; ws[1][12][4]<= -62; ws[1][12][5]<= -67; ws[1][12][6]<= 223; ws[1][12][7]<= 100; ws[1][12][8]<=-356; ws[1][12][9]<=   5; ws[1][12][10]<= 188; ws[1][12][11]<=-148; ws[1][12][12]<= 145; ws[1][12][13]<=-146; ws[1][12][14]<= -39; ws[1][12][15]<= 190;
        ws[1][13][0]<= -85; ws[1][13][1]<= 335; ws[1][13][2]<= -19; ws[1][13][3]<= -54; ws[1][13][4]<= -25; ws[1][13][5]<= 110; ws[1][13][6]<=  39; ws[1][13][7]<=-381; ws[1][13][8]<=-132; ws[1][13][9]<= -77; ws[1][13][10]<= -37; ws[1][13][11]<=-176; ws[1][13][12]<=-120; ws[1][13][13]<= 258; ws[1][13][14]<= 299; ws[1][13][15]<= 321;
        ws[1][14][0]<= 165; ws[1][14][1]<= 307; ws[1][14][2]<=-127; ws[1][14][3]<= 229; ws[1][14][4]<=  -9; ws[1][14][5]<=  70; ws[1][14][6]<= 167; ws[1][14][7]<= -80; ws[1][14][8]<= 176; ws[1][14][9]<=  21; ws[1][14][10]<=  42; ws[1][14][11]<= 271; ws[1][14][12]<= -48; ws[1][14][13]<= 228; ws[1][14][14]<=  10; ws[1][14][15]<=  10;
        ws[1][15][0]<=   3; ws[1][15][1]<=-114; ws[1][15][2]<=-301; ws[1][15][3]<= 219; ws[1][15][4]<= 172; ws[1][15][5]<= -18; ws[1][15][6]<= 376; ws[1][15][7]<=  64; ws[1][15][8]<=-193; ws[1][15][9]<=  60; ws[1][15][10]<= 249; ws[1][15][11]<=-406; ws[1][15][12]<= 260; ws[1][15][13]<= 341; ws[1][15][14]<= -73; ws[1][15][15]<=-201;

        ws[2][0 ][0]<=-173; ws[2][0 ][1]<= -25; ws[2][0 ][2]<=-142; ws[2][0 ][3]<=  97; ws[2][0 ][4]<=-150; ws[2][0 ][5]<=  17; ws[2][0 ][6]<= 457; ws[2][0 ][7]<=-345; ws[2][0 ][8]<= 250; ws[2][0 ][9]<=  -1; ws[2][0 ][10]<= 184; ws[2][0 ][11]<=  60; ws[2][0 ][12]<= 117; ws[2][0 ][13]<= 111; ws[2][0 ][14]<= -20; ws[2][0 ][15]<=-205;
        ws[2][1 ][0]<=  44; ws[2][1 ][1]<= -29; ws[2][1 ][2]<= 125; ws[2][1 ][3]<=-176; ws[2][1 ][4]<=-230; ws[2][1 ][5]<= 109; ws[2][1 ][6]<=  51; ws[2][1 ][7]<= 260; ws[2][1 ][8]<=  -3; ws[2][1 ][9]<= 120; ws[2][1 ][10]<=  26; ws[2][1 ][11]<=  -7; ws[2][1 ][12]<= 305; ws[2][1 ][13]<= 557; ws[2][1 ][14]<=  24; ws[2][1 ][15]<=  -5;
        ws[2][2 ][0]<= 214; ws[2][2 ][1]<= 107; ws[2][2 ][2]<=  91; ws[2][2 ][3]<=   8; ws[2][2 ][4]<= 263; ws[2][2 ][5]<= 130; ws[2][2 ][6]<=  29; ws[2][2 ][7]<=  -7; ws[2][2 ][8]<=  82; ws[2][2 ][9]<=   1; ws[2][2 ][10]<= 175; ws[2][2 ][11]<=  89; ws[2][2 ][12]<= 351; ws[2][2 ][13]<=-413; ws[2][2 ][14]<=  86; ws[2][2 ][15]<=-198;
        ws[2][3 ][0]<=-213; ws[2][3 ][1]<=-265; ws[2][3 ][2]<= -77; ws[2][3 ][3]<= 318; ws[2][3 ][4]<=-193; ws[2][3 ][5]<= -23; ws[2][3 ][6]<=  38; ws[2][3 ][7]<= 155; ws[2][3 ][8]<= 336; ws[2][3 ][9]<=  18; ws[2][3 ][10]<= 138; ws[2][3 ][11]<=  21; ws[2][3 ][12]<=-143; ws[2][3 ][13]<=  17; ws[2][3 ][14]<=  95; ws[2][3 ][15]<=-283;
        ws[2][4 ][0]<= 104; ws[2][4 ][1]<= 163; ws[2][4 ][2]<=-125; ws[2][4 ][3]<= -54; ws[2][4 ][4]<=-115; ws[2][4 ][5]<= 409; ws[2][4 ][6]<=  73; ws[2][4 ][7]<=  83; ws[2][4 ][8]<= -17; ws[2][4 ][9]<= 174; ws[2][4 ][10]<= 118; ws[2][4 ][11]<=-301; ws[2][4 ][12]<= -13; ws[2][4 ][13]<= 101; ws[2][4 ][14]<=-106; ws[2][4 ][15]<=  97;
        ws[2][5 ][0]<= 151; ws[2][5 ][1]<=  77; ws[2][5 ][2]<=  85; ws[2][5 ][3]<= 137; ws[2][5 ][4]<= 302; ws[2][5 ][5]<=  -5; ws[2][5 ][6]<=  93; ws[2][5 ][7]<= 235; ws[2][5 ][8]<= -19; ws[2][5 ][9]<= -59; ws[2][5 ][10]<=  14; ws[2][5 ][11]<=  44; ws[2][5 ][12]<= -97; ws[2][5 ][13]<= 192; ws[2][5 ][14]<=-357; ws[2][5 ][15]<=  -7;
        ws[2][6 ][0]<=-244; ws[2][6 ][1]<=  72; ws[2][6 ][2]<= 152; ws[2][6 ][3]<= -80; ws[2][6 ][4]<= -68; ws[2][6 ][5]<=-263; ws[2][6 ][6]<=-241; ws[2][6 ][7]<=-191; ws[2][6 ][8]<=-168; ws[2][6 ][9]<=-219; ws[2][6 ][10]<=-304; ws[2][6 ][11]<=-128; ws[2][6 ][12]<= 156; ws[2][6 ][13]<=-251; ws[2][6 ][14]<= 161; ws[2][6 ][15]<= -97;
        ws[2][7 ][0]<= -50; ws[2][7 ][1]<= -41; ws[2][7 ][2]<=-397; ws[2][7 ][3]<= -25; ws[2][7 ][4]<= -88; ws[2][7 ][5]<=  24; ws[2][7 ][6]<= 157; ws[2][7 ][7]<=-141; ws[2][7 ][8]<= 181; ws[2][7 ][9]<=-163; ws[2][7 ][10]<=  41; ws[2][7 ][11]<= 211; ws[2][7 ][12]<=-156; ws[2][7 ][13]<= -33; ws[2][7 ][14]<= 365; ws[2][7 ][15]<=-331;
        ws[2][8 ][0]<= 186; ws[2][8 ][1]<=-447; ws[2][8 ][2]<=-123; ws[2][8 ][3]<=  65; ws[2][8 ][4]<= 160; ws[2][8 ][5]<=   6; ws[2][8 ][6]<= -16; ws[2][8 ][7]<=  92; ws[2][8 ][8]<=-314; ws[2][8 ][9]<=-205; ws[2][8 ][10]<=  93; ws[2][8 ][11]<= -72; ws[2][8 ][12]<=  93; ws[2][8 ][13]<=-106; ws[2][8 ][14]<=-234; ws[2][8 ][15]<= -88;
        ws[2][9 ][0]<=  10; ws[2][9 ][1]<=-208; ws[2][9 ][2]<=   0; ws[2][9 ][3]<= -14; ws[2][9 ][4]<=  15; ws[2][9 ][5]<=-163; ws[2][9 ][6]<= -71; ws[2][9 ][7]<=  37; ws[2][9 ][8]<=  96; ws[2][9 ][9]<=  67; ws[2][9 ][10]<=-160; ws[2][9 ][11]<= 330; ws[2][9 ][12]<=  14; ws[2][9 ][13]<= 250; ws[2][9 ][14]<=-162; ws[2][9 ][15]<= 136;
        ws[2][10][0]<=-189; ws[2][10][1]<= 142; ws[2][10][2]<=-155; ws[2][10][3]<= 181; ws[2][10][4]<= 102; ws[2][10][5]<= -72; ws[2][10][6]<= 139; ws[2][10][7]<= -23; ws[2][10][8]<=  97; ws[2][10][9]<=-250; ws[2][10][10]<= 370; ws[2][10][11]<= -87; ws[2][10][12]<=  57; ws[2][10][13]<= -93; ws[2][10][14]<= -73; ws[2][10][15]<= -86;
        ws[2][11][0]<=  44; ws[2][11][1]<= 107; ws[2][11][2]<=-135; ws[2][11][3]<= -73; ws[2][11][4]<= 156; ws[2][11][5]<= 142; ws[2][11][6]<= -92; ws[2][11][7]<=  16; ws[2][11][8]<=  48; ws[2][11][9]<=-191; ws[2][11][10]<=-165; ws[2][11][11]<=  52; ws[2][11][12]<= 195; ws[2][11][13]<= 377; ws[2][11][14]<= -85; ws[2][11][15]<= 107;
        ws[2][12][0]<= -73; ws[2][12][1]<=  80; ws[2][12][2]<=  98; ws[2][12][3]<= 143; ws[2][12][4]<= -65; ws[2][12][5]<= 136; ws[2][12][6]<= 310; ws[2][12][7]<=-186; ws[2][12][8]<= 184; ws[2][12][9]<=-210; ws[2][12][10]<=-141; ws[2][12][11]<= -15; ws[2][12][12]<= 161; ws[2][12][13]<=  33; ws[2][12][14]<=-119; ws[2][12][15]<= 303;
        ws[2][13][0]<=-221; ws[2][13][1]<= -71; ws[2][13][2]<= 137; ws[2][13][3]<=-369; ws[2][13][4]<= 105; ws[2][13][5]<=  59; ws[2][13][6]<= -29; ws[2][13][7]<= -10; ws[2][13][8]<= 137; ws[2][13][9]<=-199; ws[2][13][10]<= -73; ws[2][13][11]<= -41; ws[2][13][12]<=-173; ws[2][13][13]<=-140; ws[2][13][14]<=  -6; ws[2][13][15]<=-195;
        ws[2][14][0]<= -68; ws[2][14][1]<=-187; ws[2][14][2]<= 261; ws[2][14][3]<= -72; ws[2][14][4]<= 106; ws[2][14][5]<= 164; ws[2][14][6]<= 222; ws[2][14][7]<=-192; ws[2][14][8]<=  86; ws[2][14][9]<= 175; ws[2][14][10]<= 194; ws[2][14][11]<= -91; ws[2][14][12]<= 112; ws[2][14][13]<=-141; ws[2][14][14]<= 136; ws[2][14][15]<=-140;
        ws[2][15][0]<= 153; ws[2][15][1]<=-225; ws[2][15][2]<=-115; ws[2][15][3]<=-273; ws[2][15][4]<=   8; ws[2][15][5]<=  77; ws[2][15][6]<=  32; ws[2][15][7]<= 156; ws[2][15][8]<=-123; ws[2][15][9]<= 377; ws[2][15][10]<=  12; ws[2][15][11]<=-197; ws[2][15][12]<= -63; ws[2][15][13]<= -43; ws[2][15][14]<= 219; ws[2][15][15]<= 146;

        ws[3][0 ][0]<= 302; ws[3][0 ][1]<= 136; ws[3][0 ][2]<= 122; ws[3][0 ][3]<=  56; ws[3][0 ][4]<=  41; ws[3][0 ][5]<= -87; ws[3][0 ][6]<=-310; ws[3][0 ][7]<= 240; ws[3][0 ][8]<=  78; ws[3][0 ][9]<= -85; ws[3][0 ][10]<=  24; ws[3][0 ][11]<= 284; ws[3][0 ][12]<= -41; ws[3][0 ][13]<=  13; ws[3][0 ][14]<= -48; ws[3][0 ][15]<=-218;
        ws[3][1 ][0]<= -22; ws[3][1 ][1]<=  85; ws[3][1 ][2]<=   1; ws[3][1 ][3]<= -91; ws[3][1 ][4]<= -89; ws[3][1 ][5]<=  17; ws[3][1 ][6]<= 176; ws[3][1 ][7]<= 189; ws[3][1 ][8]<=  46; ws[3][1 ][9]<= 182; ws[3][1 ][10]<=-120; ws[3][1 ][11]<=  65; ws[3][1 ][12]<= 157; ws[3][1 ][13]<= -23; ws[3][1 ][14]<=-168; ws[3][1 ][15]<=-112;
        ws[3][2 ][0]<=-147; ws[3][2 ][1]<=  36; ws[3][2 ][2]<=  19; ws[3][2 ][3]<=-182; ws[3][2 ][4]<= 101; ws[3][2 ][5]<=-225; ws[3][2 ][6]<=  88; ws[3][2 ][7]<= 217; ws[3][2 ][8]<=-186; ws[3][2 ][9]<= 129; ws[3][2 ][10]<= -43; ws[3][2 ][11]<=  63; ws[3][2 ][12]<=  67; ws[3][2 ][13]<=  13; ws[3][2 ][14]<= 196; ws[3][2 ][15]<=-237;
        ws[3][3 ][0]<=-125; ws[3][3 ][1]<= 282; ws[3][3 ][2]<= 133; ws[3][3 ][3]<= 160; ws[3][3 ][4]<=-312; ws[3][3 ][5]<=   4; ws[3][3 ][6]<=-146; ws[3][3 ][7]<=  70; ws[3][3 ][8]<= 120; ws[3][3 ][9]<=-173; ws[3][3 ][10]<= 172; ws[3][3 ][11]<= 189; ws[3][3 ][12]<=   1; ws[3][3 ][13]<=-141; ws[3][3 ][14]<= -59; ws[3][3 ][15]<=  74;
        ws[3][4 ][0]<=  13; ws[3][4 ][1]<=  91; ws[3][4 ][2]<= 114; ws[3][4 ][3]<= 196; ws[3][4 ][4]<= 170; ws[3][4 ][5]<= -66; ws[3][4 ][6]<=-213; ws[3][4 ][7]<= -91; ws[3][4 ][8]<=-199; ws[3][4 ][9]<=-274; ws[3][4 ][10]<=-296; ws[3][4 ][11]<=  94; ws[3][4 ][12]<=-257; ws[3][4 ][13]<=-161; ws[3][4 ][14]<= 190; ws[3][4 ][15]<= -30;
        ws[3][5 ][0]<= 388; ws[3][5 ][1]<= 260; ws[3][5 ][2]<=  85; ws[3][5 ][3]<=-326; ws[3][5 ][4]<=  -8; ws[3][5 ][5]<=  62; ws[3][5 ][6]<= 160; ws[3][5 ][7]<=-111; ws[3][5 ][8]<= 260; ws[3][5 ][9]<=-216; ws[3][5 ][10]<= -98; ws[3][5 ][11]<= -13; ws[3][5 ][12]<= -34; ws[3][5 ][13]<=-160; ws[3][5 ][14]<= 178; ws[3][5 ][15]<= -20;
        ws[3][6 ][0]<=-264; ws[3][6 ][1]<= 130; ws[3][6 ][2]<= -71; ws[3][6 ][3]<=  67; ws[3][6 ][4]<=-189; ws[3][6 ][5]<=  78; ws[3][6 ][6]<= 141; ws[3][6 ][7]<= 234; ws[3][6 ][8]<=-230; ws[3][6 ][9]<=-210; ws[3][6 ][10]<= -59; ws[3][6 ][11]<= 169; ws[3][6 ][12]<= -61; ws[3][6 ][13]<=-165; ws[3][6 ][14]<= 138; ws[3][6 ][15]<=-238;
        ws[3][7 ][0]<= -78; ws[3][7 ][1]<=  63; ws[3][7 ][2]<= -88; ws[3][7 ][3]<= 333; ws[3][7 ][4]<=  86; ws[3][7 ][5]<= -34; ws[3][7 ][6]<=  39; ws[3][7 ][7]<= -86; ws[3][7 ][8]<=-185; ws[3][7 ][9]<=-112; ws[3][7 ][10]<= 286; ws[3][7 ][11]<=-362; ws[3][7 ][12]<= 158; ws[3][7 ][13]<=  72; ws[3][7 ][14]<= -65; ws[3][7 ][15]<=  88;
        ws[3][8 ][0]<= -31; ws[3][8 ][1]<=-202; ws[3][8 ][2]<= 185; ws[3][8 ][3]<=-184; ws[3][8 ][4]<=-120; ws[3][8 ][5]<= 336; ws[3][8 ][6]<= -21; ws[3][8 ][7]<= 143; ws[3][8 ][8]<= 233; ws[3][8 ][9]<=  -9; ws[3][8 ][10]<= 144; ws[3][8 ][11]<=  63; ws[3][8 ][12]<= -38; ws[3][8 ][13]<= 332; ws[3][8 ][14]<= -77; ws[3][8 ][15]<= 329;
        ws[3][9 ][0]<= -74; ws[3][9 ][1]<=  48; ws[3][9 ][2]<=-300; ws[3][9 ][3]<= -73; ws[3][9 ][4]<=-295; ws[3][9 ][5]<=-372; ws[3][9 ][6]<= -34; ws[3][9 ][7]<=   5; ws[3][9 ][8]<= 159; ws[3][9 ][9]<= 106; ws[3][9 ][10]<=-121; ws[3][9 ][11]<= -68; ws[3][9 ][12]<=-102; ws[3][9 ][13]<= 214; ws[3][9 ][14]<= -52; ws[3][9 ][15]<= 139;
        ws[3][10][0]<=-176; ws[3][10][1]<= -72; ws[3][10][2]<= 144; ws[3][10][3]<=  55; ws[3][10][4]<= -50; ws[3][10][5]<=-294; ws[3][10][6]<=  19; ws[3][10][7]<=-154; ws[3][10][8]<= 169; ws[3][10][9]<= 262; ws[3][10][10]<=  21; ws[3][10][11]<= 221; ws[3][10][12]<= 171; ws[3][10][13]<= 375; ws[3][10][14]<= 244; ws[3][10][15]<=  99;
        ws[3][11][0]<=  -8; ws[3][11][1]<=   3; ws[3][11][2]<=  -9; ws[3][11][3]<= 265; ws[3][11][4]<=  70; ws[3][11][5]<= 207; ws[3][11][6]<=   7; ws[3][11][7]<=  38; ws[3][11][8]<= -12; ws[3][11][9]<=-204; ws[3][11][10]<=-124; ws[3][11][11]<=-140; ws[3][11][12]<= 297; ws[3][11][13]<= 130; ws[3][11][14]<=   6; ws[3][11][15]<=-138;
        ws[3][12][0]<= 146; ws[3][12][1]<=-145; ws[3][12][2]<= 192; ws[3][12][3]<=  36; ws[3][12][4]<= 270; ws[3][12][5]<= 197; ws[3][12][6]<= 182; ws[3][12][7]<=  20; ws[3][12][8]<=-188; ws[3][12][9]<= -82; ws[3][12][10]<=-242; ws[3][12][11]<= 300; ws[3][12][12]<=-310; ws[3][12][13]<=  12; ws[3][12][14]<=  21; ws[3][12][15]<= -97;
        ws[3][13][0]<=-109; ws[3][13][1]<= 138; ws[3][13][2]<=  89; ws[3][13][3]<= -24; ws[3][13][4]<= -47; ws[3][13][5]<=  12; ws[3][13][6]<=-208; ws[3][13][7]<=-299; ws[3][13][8]<= -78; ws[3][13][9]<= -39; ws[3][13][10]<=  76; ws[3][13][11]<= -43; ws[3][13][12]<= 372; ws[3][13][13]<= -86; ws[3][13][14]<= 112; ws[3][13][15]<=-220;
        ws[3][14][0]<= 322; ws[3][14][1]<=-219; ws[3][14][2]<=-169; ws[3][14][3]<= 181; ws[3][14][4]<= 156; ws[3][14][5]<= 184; ws[3][14][6]<= -93; ws[3][14][7]<=-148; ws[3][14][8]<= -23; ws[3][14][9]<=  52; ws[3][14][10]<= 130; ws[3][14][11]<=  37; ws[3][14][12]<= 108; ws[3][14][13]<= 167; ws[3][14][14]<= 235; ws[3][14][15]<= -50;
        ws[3][15][0]<=  10; ws[3][15][1]<=-271; ws[3][15][2]<=-386; ws[3][15][3]<=-153; ws[3][15][4]<= -54; ws[3][15][5]<=  17; ws[3][15][6]<=-118; ws[3][15][7]<=   9; ws[3][15][8]<= 148; ws[3][15][9]<= 112; ws[3][15][10]<=-121; ws[3][15][11]<=-164; ws[3][15][12]<=  84; ws[3][15][13]<=-176; ws[3][15][14]<=  41; ws[3][15][15]<= 224;

        ws[4][0 ][0]<= -21; ws[4][0 ][1]<= 130; ws[4][0 ][2]<= 176; ws[4][0 ][3]<= -31; ws[4][0 ][4]<=  28; ws[4][0 ][5]<=-115; ws[4][0 ][6]<= 256; ws[4][0 ][7]<=  44; ws[4][0 ][8]<=-313; ws[4][0 ][9]<= 258; ws[4][0 ][10]<= 193; ws[4][0 ][11]<= -91; ws[4][0 ][12]<= -17; ws[4][0 ][13]<= 172; ws[4][0 ][14]<=  50; ws[4][0 ][15]<= 167;
        ws[4][1 ][0]<= -31; ws[4][1 ][1]<= -89; ws[4][1 ][2]<= -84; ws[4][1 ][3]<=-168; ws[4][1 ][4]<=  23; ws[4][1 ][5]<=-407; ws[4][1 ][6]<= -14; ws[4][1 ][7]<= 105; ws[4][1 ][8]<=  22; ws[4][1 ][9]<=-101; ws[4][1 ][10]<=  68; ws[4][1 ][11]<= -64; ws[4][1 ][12]<=-485; ws[4][1 ][13]<=-391; ws[4][1 ][14]<=  94; ws[4][1 ][15]<=-210;
        ws[4][2 ][0]<=-385; ws[4][2 ][1]<= 360; ws[4][2 ][2]<=-199; ws[4][2 ][3]<=-222; ws[4][2 ][4]<=-256; ws[4][2 ][5]<= 171; ws[4][2 ][6]<=-179; ws[4][2 ][7]<=  83; ws[4][2 ][8]<= -54; ws[4][2 ][9]<= 197; ws[4][2 ][10]<= 188; ws[4][2 ][11]<=-282; ws[4][2 ][12]<= -29; ws[4][2 ][13]<= 300; ws[4][2 ][14]<=-124; ws[4][2 ][15]<= 217;
        ws[4][3 ][0]<=  57; ws[4][3 ][1]<=  17; ws[4][3 ][2]<=-195; ws[4][3 ][3]<= 177; ws[4][3 ][4]<= 147; ws[4][3 ][5]<=-128; ws[4][3 ][6]<= -10; ws[4][3 ][7]<= 172; ws[4][3 ][8]<= -75; ws[4][3 ][9]<= 202; ws[4][3 ][10]<= -64; ws[4][3 ][11]<= -76; ws[4][3 ][12]<=-310; ws[4][3 ][13]<= 139; ws[4][3 ][14]<= -37; ws[4][3 ][15]<=-158;
        ws[4][4 ][0]<= 179; ws[4][4 ][1]<= 205; ws[4][4 ][2]<= 258; ws[4][4 ][3]<= 319; ws[4][4 ][4]<=  26; ws[4][4 ][5]<= 160; ws[4][4 ][6]<=-273; ws[4][4 ][7]<= -10; ws[4][4 ][8]<= 113; ws[4][4 ][9]<= 213; ws[4][4 ][10]<= 167; ws[4][4 ][11]<=-494; ws[4][4 ][12]<=  98; ws[4][4 ][13]<= 299; ws[4][4 ][14]<=-288; ws[4][4 ][15]<=-208;
        ws[4][5 ][0]<=-112; ws[4][5 ][1]<=  11; ws[4][5 ][2]<= -98; ws[4][5 ][3]<=  33; ws[4][5 ][4]<=  82; ws[4][5 ][5]<=-459; ws[4][5 ][6]<=-164; ws[4][5 ][7]<=-202; ws[4][5 ][8]<= -16; ws[4][5 ][9]<=-433; ws[4][5 ][10]<=-262; ws[4][5 ][11]<=   1; ws[4][5 ][12]<=-228; ws[4][5 ][13]<= 127; ws[4][5 ][14]<=-159; ws[4][5 ][15]<=-157;
        ws[4][6 ][0]<=-191; ws[4][6 ][1]<=-148; ws[4][6 ][2]<=  52; ws[4][6 ][3]<=  70; ws[4][6 ][4]<= -93; ws[4][6 ][5]<= -93; ws[4][6 ][6]<=-291; ws[4][6 ][7]<=  53; ws[4][6 ][8]<=-239; ws[4][6 ][9]<=-151; ws[4][6 ][10]<=  50; ws[4][6 ][11]<= 224; ws[4][6 ][12]<=  13; ws[4][6 ][13]<= -28; ws[4][6 ][14]<=-120; ws[4][6 ][15]<=  90;
        ws[4][7 ][0]<=-176; ws[4][7 ][1]<=-201; ws[4][7 ][2]<= -54; ws[4][7 ][3]<=-242; ws[4][7 ][4]<= 189; ws[4][7 ][5]<=-142; ws[4][7 ][6]<= -58; ws[4][7 ][7]<= -74; ws[4][7 ][8]<=-261; ws[4][7 ][9]<=   9; ws[4][7 ][10]<=-206; ws[4][7 ][11]<=  -9; ws[4][7 ][12]<=  23; ws[4][7 ][13]<=  -2; ws[4][7 ][14]<=-279; ws[4][7 ][15]<=  85;
        ws[4][8 ][0]<=-170; ws[4][8 ][1]<=  21; ws[4][8 ][2]<=   2; ws[4][8 ][3]<= -79; ws[4][8 ][4]<= 196; ws[4][8 ][5]<= -57; ws[4][8 ][6]<=  13; ws[4][8 ][7]<= 179; ws[4][8 ][8]<= 237; ws[4][8 ][9]<= -53; ws[4][8 ][10]<=-147; ws[4][8 ][11]<= 244; ws[4][8 ][12]<= 176; ws[4][8 ][13]<=  97; ws[4][8 ][14]<=-100; ws[4][8 ][15]<=  12;
        ws[4][9 ][0]<=  99; ws[4][9 ][1]<=-104; ws[4][9 ][2]<=  94; ws[4][9 ][3]<= -77; ws[4][9 ][4]<= 138; ws[4][9 ][5]<=  86; ws[4][9 ][6]<= -35; ws[4][9 ][7]<=-149; ws[4][9 ][8]<=-139; ws[4][9 ][9]<= -84; ws[4][9 ][10]<=  20; ws[4][9 ][11]<= -54; ws[4][9 ][12]<= 193; ws[4][9 ][13]<=  14; ws[4][9 ][14]<=-130; ws[4][9 ][15]<= -94;
        ws[4][10][0]<=-202; ws[4][10][1]<= 178; ws[4][10][2]<=  21; ws[4][10][3]<=-170; ws[4][10][4]<=-209; ws[4][10][5]<= -79; ws[4][10][6]<= -45; ws[4][10][7]<= 108; ws[4][10][8]<=   4; ws[4][10][9]<=   3; ws[4][10][10]<=-179; ws[4][10][11]<=  60; ws[4][10][12]<=  90; ws[4][10][13]<= 197; ws[4][10][14]<= 204; ws[4][10][15]<= 240;
        ws[4][11][0]<= -26; ws[4][11][1]<=-125; ws[4][11][2]<= -17; ws[4][11][3]<=-131; ws[4][11][4]<= 195; ws[4][11][5]<= -57; ws[4][11][6]<= 189; ws[4][11][7]<=-203; ws[4][11][8]<= 156; ws[4][11][9]<= 169; ws[4][11][10]<=-105; ws[4][11][11]<=-197; ws[4][11][12]<=  75; ws[4][11][13]<= 220; ws[4][11][14]<=  45; ws[4][11][15]<=   5;
        ws[4][12][0]<= 152; ws[4][12][1]<=  93; ws[4][12][2]<=-304; ws[4][12][3]<= -31; ws[4][12][4]<= 292; ws[4][12][5]<= -88; ws[4][12][6]<= -30; ws[4][12][7]<=  65; ws[4][12][8]<= 160; ws[4][12][9]<=-161; ws[4][12][10]<= 233; ws[4][12][11]<=   5; ws[4][12][12]<=  62; ws[4][12][13]<=  99; ws[4][12][14]<= -36; ws[4][12][15]<=-266;
        ws[4][13][0]<= 150; ws[4][13][1]<= 104; ws[4][13][2]<= 155; ws[4][13][3]<=   6; ws[4][13][4]<= -60; ws[4][13][5]<=-283; ws[4][13][6]<=-276; ws[4][13][7]<= 397; ws[4][13][8]<= 177; ws[4][13][9]<=  -8; ws[4][13][10]<= -77; ws[4][13][11]<= -21; ws[4][13][12]<=   0; ws[4][13][13]<=  35; ws[4][13][14]<= 232; ws[4][13][15]<=  25;
        ws[4][14][0]<=  82; ws[4][14][1]<= -51; ws[4][14][2]<= 252; ws[4][14][3]<= -46; ws[4][14][4]<=-185; ws[4][14][5]<=  79; ws[4][14][6]<=  94; ws[4][14][7]<=-181; ws[4][14][8]<= 264; ws[4][14][9]<= -89; ws[4][14][10]<= -54; ws[4][14][11]<=-199; ws[4][14][12]<=  64; ws[4][14][13]<=  68; ws[4][14][14]<=  69; ws[4][14][15]<= 126;
        ws[4][15][0]<=  39; ws[4][15][1]<= 302; ws[4][15][2]<=  53; ws[4][15][3]<=-170; ws[4][15][4]<= -83; ws[4][15][5]<= -59; ws[4][15][6]<=  64; ws[4][15][7]<=-210; ws[4][15][8]<=  81; ws[4][15][9]<= 234; ws[4][15][10]<= 200; ws[4][15][11]<=-258; ws[4][15][12]<= 113; ws[4][15][13]<=  -9; ws[4][15][14]<=-206; ws[4][15][15]<=-134;

        ws[5][0 ][0]<= 157; ws[5][0 ][1]<=-152; ws[5][0 ][2]<= -36; ws[5][0 ][3]<=-198; ws[5][0 ][4]<= 322; ws[5][0 ][5]<= 271; ws[5][0 ][6]<=-375; ws[5][0 ][7]<=-109; ws[5][0 ][8]<= 368; ws[5][0 ][9]<=-122; ws[5][0 ][10]<=  65; ws[5][0 ][11]<=  55; ws[5][0 ][12]<=-244; ws[5][0 ][13]<=  14; ws[5][0 ][14]<=  87; ws[5][0 ][15]<=-136;
        ws[5][1 ][0]<=  55; ws[5][1 ][1]<=  61; ws[5][1 ][2]<= 243; ws[5][1 ][3]<=   0; ws[5][1 ][4]<=  41; ws[5][1 ][5]<=  87; ws[5][1 ][6]<=  92; ws[5][1 ][7]<= 146; ws[5][1 ][8]<=   3; ws[5][1 ][9]<= 131; ws[5][1 ][10]<=  -1; ws[5][1 ][11]<= 152; ws[5][1 ][12]<=-239; ws[5][1 ][13]<= -44; ws[5][1 ][14]<= 384; ws[5][1 ][15]<= 235;
        ws[5][2 ][0]<= 142; ws[5][2 ][1]<=  75; ws[5][2 ][2]<= -33; ws[5][2 ][3]<=  77; ws[5][2 ][4]<= -72; ws[5][2 ][5]<= 271; ws[5][2 ][6]<=-199; ws[5][2 ][7]<=   8; ws[5][2 ][8]<= 174; ws[5][2 ][9]<=-100; ws[5][2 ][10]<= 202; ws[5][2 ][11]<=-119; ws[5][2 ][12]<= 129; ws[5][2 ][13]<=  67; ws[5][2 ][14]<=-229; ws[5][2 ][15]<= -43;
        ws[5][3 ][0]<= -79; ws[5][3 ][1]<= -49; ws[5][3 ][2]<= -18; ws[5][3 ][3]<= -37; ws[5][3 ][4]<=  38; ws[5][3 ][5]<=  -1; ws[5][3 ][6]<=-126; ws[5][3 ][7]<= 194; ws[5][3 ][8]<=  23; ws[5][3 ][9]<=-238; ws[5][3 ][10]<=   6; ws[5][3 ][11]<= -53; ws[5][3 ][12]<= 188; ws[5][3 ][13]<=-198; ws[5][3 ][14]<=-111; ws[5][3 ][15]<=-148;
        ws[5][4 ][0]<= 166; ws[5][4 ][1]<= 115; ws[5][4 ][2]<=-227; ws[5][4 ][3]<=  84; ws[5][4 ][4]<=-144; ws[5][4 ][5]<=-146; ws[5][4 ][6]<= -44; ws[5][4 ][7]<=-190; ws[5][4 ][8]<=-347; ws[5][4 ][9]<=  91; ws[5][4 ][10]<=  67; ws[5][4 ][11]<=-178; ws[5][4 ][12]<= 121; ws[5][4 ][13]<=-118; ws[5][4 ][14]<=  11; ws[5][4 ][15]<=-109;
        ws[5][5 ][0]<=-383; ws[5][5 ][1]<=  17; ws[5][5 ][2]<=-130; ws[5][5 ][3]<=-137; ws[5][5 ][4]<=-116; ws[5][5 ][5]<= 130; ws[5][5 ][6]<=-108; ws[5][5 ][7]<= -48; ws[5][5 ][8]<=  20; ws[5][5 ][9]<= 206; ws[5][5 ][10]<=-105; ws[5][5 ][11]<=-108; ws[5][5 ][12]<=  40; ws[5][5 ][13]<=-169; ws[5][5 ][14]<= -36; ws[5][5 ][15]<= -38;
        ws[5][6 ][0]<=  76; ws[5][6 ][1]<=-164; ws[5][6 ][2]<=-109; ws[5][6 ][3]<= 282; ws[5][6 ][4]<=-221; ws[5][6 ][5]<=  21; ws[5][6 ][6]<= -71; ws[5][6 ][7]<=-125; ws[5][6 ][8]<= 231; ws[5][6 ][9]<=-120; ws[5][6 ][10]<= -64; ws[5][6 ][11]<=-173; ws[5][6 ][12]<= 380; ws[5][6 ][13]<=-377; ws[5][6 ][14]<=   6; ws[5][6 ][15]<=-278;
        ws[5][7 ][0]<= -38; ws[5][7 ][1]<= 149; ws[5][7 ][2]<=  49; ws[5][7 ][3]<= 152; ws[5][7 ][4]<= -26; ws[5][7 ][5]<= -54; ws[5][7 ][6]<=-138; ws[5][7 ][7]<= -72; ws[5][7 ][8]<=-111; ws[5][7 ][9]<=-157; ws[5][7 ][10]<= 393; ws[5][7 ][11]<= 228; ws[5][7 ][12]<= 116; ws[5][7 ][13]<= 145; ws[5][7 ][14]<= 194; ws[5][7 ][15]<= -98;
        ws[5][8 ][0]<= -55; ws[5][8 ][1]<= 252; ws[5][8 ][2]<= -10; ws[5][8 ][3]<= -19; ws[5][8 ][4]<= 361; ws[5][8 ][5]<= 243; ws[5][8 ][6]<=  54; ws[5][8 ][7]<= -65; ws[5][8 ][8]<=-136; ws[5][8 ][9]<=-166; ws[5][8 ][10]<= 155; ws[5][8 ][11]<=  37; ws[5][8 ][12]<= -49; ws[5][8 ][13]<=-348; ws[5][8 ][14]<= 194; ws[5][8 ][15]<= 193;
        ws[5][9 ][0]<=  -8; ws[5][9 ][1]<= 211; ws[5][9 ][2]<=-359; ws[5][9 ][3]<= 170; ws[5][9 ][4]<=-159; ws[5][9 ][5]<=-244; ws[5][9 ][6]<=-118; ws[5][9 ][7]<=  -2; ws[5][9 ][8]<= 175; ws[5][9 ][9]<= -80; ws[5][9 ][10]<=-237; ws[5][9 ][11]<= 345; ws[5][9 ][12]<= 189; ws[5][9 ][13]<=-149; ws[5][9 ][14]<= 147; ws[5][9 ][15]<= -50;
        ws[5][10][0]<= 132; ws[5][10][1]<= -53; ws[5][10][2]<=   2; ws[5][10][3]<=  50; ws[5][10][4]<= -21; ws[5][10][5]<= -88; ws[5][10][6]<=-117; ws[5][10][7]<=  74; ws[5][10][8]<=  55; ws[5][10][9]<=-368; ws[5][10][10]<=-348; ws[5][10][11]<= 218; ws[5][10][12]<=  96; ws[5][10][13]<= 334; ws[5][10][14]<= -15; ws[5][10][15]<= 241;
        ws[5][11][0]<=  37; ws[5][11][1]<=-177; ws[5][11][2]<=  28; ws[5][11][3]<=-374; ws[5][11][4]<= 119; ws[5][11][5]<= 132; ws[5][11][6]<=-331; ws[5][11][7]<=-443; ws[5][11][8]<= 174; ws[5][11][9]<=-263; ws[5][11][10]<=-130; ws[5][11][11]<= -66; ws[5][11][12]<= -36; ws[5][11][13]<= 128; ws[5][11][14]<=-314; ws[5][11][15]<=-237;
        ws[5][12][0]<= 182; ws[5][12][1]<= -39; ws[5][12][2]<=-241; ws[5][12][3]<=-125; ws[5][12][4]<=-315; ws[5][12][5]<= -19; ws[5][12][6]<= 184; ws[5][12][7]<=-141; ws[5][12][8]<= 177; ws[5][12][9]<= 156; ws[5][12][10]<=-234; ws[5][12][11]<=  63; ws[5][12][12]<= 156; ws[5][12][13]<=  86; ws[5][12][14]<=  84; ws[5][12][15]<=  33;
        ws[5][13][0]<=-190; ws[5][13][1]<= 190; ws[5][13][2]<=-303; ws[5][13][3]<=  10; ws[5][13][4]<= 138; ws[5][13][5]<= 167; ws[5][13][6]<=-142; ws[5][13][7]<=-141; ws[5][13][8]<=  41; ws[5][13][9]<=-162; ws[5][13][10]<=  48; ws[5][13][11]<= 275; ws[5][13][12]<=  21; ws[5][13][13]<=-361; ws[5][13][14]<=-189; ws[5][13][15]<=-189;
        ws[5][14][0]<= 132; ws[5][14][1]<=  58; ws[5][14][2]<= 276; ws[5][14][3]<= -51; ws[5][14][4]<=-259; ws[5][14][5]<=  10; ws[5][14][6]<= 134; ws[5][14][7]<= 156; ws[5][14][8]<=-404; ws[5][14][9]<= 146; ws[5][14][10]<=-133; ws[5][14][11]<= 114; ws[5][14][12]<=  -2; ws[5][14][13]<= -79; ws[5][14][14]<=-210; ws[5][14][15]<= 142;
        ws[5][15][0]<=-304; ws[5][15][1]<=-421; ws[5][15][2]<=-134; ws[5][15][3]<= 109; ws[5][15][4]<=-118; ws[5][15][5]<= 103; ws[5][15][6]<=  48; ws[5][15][7]<= -26; ws[5][15][8]<=  78; ws[5][15][9]<= -80; ws[5][15][10]<= -52; ws[5][15][11]<= -59; ws[5][15][12]<= -95; ws[5][15][13]<=  95; ws[5][15][14]<=  53; ws[5][15][15]<=-160;

        ws[6][0 ][0]<= -95; ws[6][0 ][1]<=-167; ws[6][0 ][2]<= 148; ws[6][0 ][3]<= 138; ws[6][0 ][4]<=-287; ws[6][0 ][5]<= -56; ws[6][0 ][6]<= -14; ws[6][0 ][7]<= 282; ws[6][0 ][8]<= 137; ws[6][0 ][9]<=  54; ws[6][0 ][10]<=-469; ws[6][0 ][11]<=-420; ws[6][0 ][12]<=-343; ws[6][0 ][13]<= 194; ws[6][0 ][14]<=-362; ws[6][0 ][15]<=  28;
        ws[6][1 ][0]<= -45; ws[6][1 ][1]<=  81; ws[6][1 ][2]<=  69; ws[6][1 ][3]<= 347; ws[6][1 ][4]<= -22; ws[6][1 ][5]<=  98; ws[6][1 ][6]<=  30; ws[6][1 ][7]<= 322; ws[6][1 ][8]<= -15; ws[6][1 ][9]<= -14; ws[6][1 ][10]<= 117; ws[6][1 ][11]<=   3; ws[6][1 ][12]<=  63; ws[6][1 ][13]<=  49; ws[6][1 ][14]<= 212; ws[6][1 ][15]<=-130;
        ws[6][2 ][0]<= 238; ws[6][2 ][1]<= 424; ws[6][2 ][2]<= -46; ws[6][2 ][3]<=  -2; ws[6][2 ][4]<= -69; ws[6][2 ][5]<= -22; ws[6][2 ][6]<= 224; ws[6][2 ][7]<= 132; ws[6][2 ][8]<= 133; ws[6][2 ][9]<= 354; ws[6][2 ][10]<=  21; ws[6][2 ][11]<=  28; ws[6][2 ][12]<=-144; ws[6][2 ][13]<= -44; ws[6][2 ][14]<= 123; ws[6][2 ][15]<=-211;
        ws[6][3 ][0]<=-442; ws[6][3 ][1]<=-213; ws[6][3 ][2]<=  94; ws[6][3 ][3]<= -93; ws[6][3 ][4]<=  61; ws[6][3 ][5]<= -45; ws[6][3 ][6]<=-144; ws[6][3 ][7]<=-243; ws[6][3 ][8]<=-131; ws[6][3 ][9]<= -80; ws[6][3 ][10]<=  -4; ws[6][3 ][11]<=  -2; ws[6][3 ][12]<=-332; ws[6][3 ][13]<=  37; ws[6][3 ][14]<=-153; ws[6][3 ][15]<=-424;
        ws[6][4 ][0]<=-104; ws[6][4 ][1]<=   0; ws[6][4 ][2]<= -12; ws[6][4 ][3]<= -89; ws[6][4 ][4]<=  55; ws[6][4 ][5]<= 231; ws[6][4 ][6]<= -64; ws[6][4 ][7]<=-314; ws[6][4 ][8]<= 241; ws[6][4 ][9]<= 253; ws[6][4 ][10]<=-150; ws[6][4 ][11]<= -49; ws[6][4 ][12]<= -43; ws[6][4 ][13]<=  25; ws[6][4 ][14]<= -61; ws[6][4 ][15]<= 130;
        ws[6][5 ][0]<= -14; ws[6][5 ][1]<=-280; ws[6][5 ][2]<= 146; ws[6][5 ][3]<=  68; ws[6][5 ][4]<= -94; ws[6][5 ][5]<= 196; ws[6][5 ][6]<=-122; ws[6][5 ][7]<=  56; ws[6][5 ][8]<= -99; ws[6][5 ][9]<=-149; ws[6][5 ][10]<=  52; ws[6][5 ][11]<=  53; ws[6][5 ][12]<=  24; ws[6][5 ][13]<= 182; ws[6][5 ][14]<= 164; ws[6][5 ][15]<= 220;
        ws[6][6 ][0]<=  38; ws[6][6 ][1]<= -15; ws[6][6 ][2]<=-220; ws[6][6 ][3]<=-196; ws[6][6 ][4]<=  10; ws[6][6 ][5]<= -14; ws[6][6 ][6]<=-321; ws[6][6 ][7]<= -36; ws[6][6 ][8]<=-303; ws[6][6 ][9]<=-194; ws[6][6 ][10]<=  -4; ws[6][6 ][11]<=  16; ws[6][6 ][12]<=-143; ws[6][6 ][13]<=-276; ws[6][6 ][14]<= -68; ws[6][6 ][15]<= 131;
        ws[6][7 ][0]<= -93; ws[6][7 ][1]<= -80; ws[6][7 ][2]<=  31; ws[6][7 ][3]<= -22; ws[6][7 ][4]<= -54; ws[6][7 ][5]<= 337; ws[6][7 ][6]<= 244; ws[6][7 ][7]<=  42; ws[6][7 ][8]<= -39; ws[6][7 ][9]<= -65; ws[6][7 ][10]<=  -5; ws[6][7 ][11]<= 283; ws[6][7 ][12]<= -39; ws[6][7 ][13]<= 133; ws[6][7 ][14]<= 153; ws[6][7 ][15]<= 197;
        ws[6][8 ][0]<=  99; ws[6][8 ][1]<= -50; ws[6][8 ][2]<= 280; ws[6][8 ][3]<= -14; ws[6][8 ][4]<= 273; ws[6][8 ][5]<=   5; ws[6][8 ][6]<=-229; ws[6][8 ][7]<= 108; ws[6][8 ][8]<= -84; ws[6][8 ][9]<= 110; ws[6][8 ][10]<=  30; ws[6][8 ][11]<=  28; ws[6][8 ][12]<= -49; ws[6][8 ][13]<= 323; ws[6][8 ][14]<=-112; ws[6][8 ][15]<= 269;
        ws[6][9 ][0]<= 197; ws[6][9 ][1]<= -17; ws[6][9 ][2]<=  29; ws[6][9 ][3]<= 137; ws[6][9 ][4]<=-167; ws[6][9 ][5]<= 199; ws[6][9 ][6]<= 163; ws[6][9 ][7]<=  15; ws[6][9 ][8]<= 239; ws[6][9 ][9]<= 307; ws[6][9 ][10]<= 127; ws[6][9 ][11]<=-109; ws[6][9 ][12]<=  13; ws[6][9 ][13]<= -96; ws[6][9 ][14]<= -73; ws[6][9 ][15]<= -62;
        ws[6][10][0]<= -58; ws[6][10][1]<=-240; ws[6][10][2]<=  39; ws[6][10][3]<=   9; ws[6][10][4]<= -49; ws[6][10][5]<= 240; ws[6][10][6]<= -48; ws[6][10][7]<=  38; ws[6][10][8]<=  15; ws[6][10][9]<=-202; ws[6][10][10]<= 230; ws[6][10][11]<= 247; ws[6][10][12]<= 101; ws[6][10][13]<= 179; ws[6][10][14]<= 157; ws[6][10][15]<= 169;
        ws[6][11][0]<= 120; ws[6][11][1]<=  52; ws[6][11][2]<= 234; ws[6][11][3]<= -87; ws[6][11][4]<=-205; ws[6][11][5]<=-178; ws[6][11][6]<=  94; ws[6][11][7]<= 189; ws[6][11][8]<=-123; ws[6][11][9]<=  16; ws[6][11][10]<= -30; ws[6][11][11]<=-101; ws[6][11][12]<= 142; ws[6][11][13]<= 288; ws[6][11][14]<=  40; ws[6][11][15]<=   5;
        ws[6][12][0]<=  54; ws[6][12][1]<=-117; ws[6][12][2]<= 366; ws[6][12][3]<= -32; ws[6][12][4]<=  49; ws[6][12][5]<=  50; ws[6][12][6]<= -75; ws[6][12][7]<= 400; ws[6][12][8]<= 267; ws[6][12][9]<= -43; ws[6][12][10]<= -91; ws[6][12][11]<= -41; ws[6][12][12]<= -23; ws[6][12][13]<=  94; ws[6][12][14]<= -74; ws[6][12][15]<= 252;
        ws[6][13][0]<=  75; ws[6][13][1]<=  44; ws[6][13][2]<=   5; ws[6][13][3]<=-165; ws[6][13][4]<=  66; ws[6][13][5]<=-238; ws[6][13][6]<=  74; ws[6][13][7]<= 106; ws[6][13][8]<= -29; ws[6][13][9]<= -16; ws[6][13][10]<=   2; ws[6][13][11]<=  74; ws[6][13][12]<=  66; ws[6][13][13]<= 136; ws[6][13][14]<=   3; ws[6][13][15]<=  93;
        ws[6][14][0]<=-134; ws[6][14][1]<= 177; ws[6][14][2]<= 255; ws[6][14][3]<= 279; ws[6][14][4]<=  14; ws[6][14][5]<= 278; ws[6][14][6]<= 415; ws[6][14][7]<=  -4; ws[6][14][8]<= 314; ws[6][14][9]<= 165; ws[6][14][10]<=  -7; ws[6][14][11]<=   0; ws[6][14][12]<=-139; ws[6][14][13]<= -55; ws[6][14][14]<=  -6; ws[6][14][15]<=-306;
        ws[6][15][0]<= 103; ws[6][15][1]<= -51; ws[6][15][2]<=   5; ws[6][15][3]<=  36; ws[6][15][4]<=  64; ws[6][15][5]<=-121; ws[6][15][6]<=   8; ws[6][15][7]<=  48; ws[6][15][8]<=  55; ws[6][15][9]<= 328; ws[6][15][10]<= -49; ws[6][15][11]<= -47; ws[6][15][12]<= -51; ws[6][15][13]<=-225; ws[6][15][14]<=-125; ws[6][15][15]<= 280;

        ws[7][0 ][0]<= 236; ws[7][0 ][1]<=-127; ws[7][0 ][2]<=-339; ws[7][0 ][3]<= 149; ws[7][0 ][4]<=   5; ws[7][0 ][5]<=-341; ws[7][0 ][6]<= -60; ws[7][0 ][7]<=  22; ws[7][0 ][8]<= -56; ws[7][0 ][9]<=-233; ws[7][0 ][10]<= 117; ws[7][0 ][11]<= 122; ws[7][0 ][12]<=  23; ws[7][0 ][13]<=-172; ws[7][0 ][14]<= 181; ws[7][0 ][15]<=-109;
        ws[7][1 ][0]<=  23; ws[7][1 ][1]<= -78; ws[7][1 ][2]<=  74; ws[7][1 ][3]<=-197; ws[7][1 ][4]<=-142; ws[7][1 ][5]<= 142; ws[7][1 ][6]<=  19; ws[7][1 ][7]<= -34; ws[7][1 ][8]<=-367; ws[7][1 ][9]<=  37; ws[7][1 ][10]<= 123; ws[7][1 ][11]<=-100; ws[7][1 ][12]<= -67; ws[7][1 ][13]<=-297; ws[7][1 ][14]<=  -4; ws[7][1 ][15]<=  -9;
        ws[7][2 ][0]<=  81; ws[7][2 ][1]<= -77; ws[7][2 ][2]<=-206; ws[7][2 ][3]<= -19; ws[7][2 ][4]<=-242; ws[7][2 ][5]<= -49; ws[7][2 ][6]<= 184; ws[7][2 ][7]<=  13; ws[7][2 ][8]<= 236; ws[7][2 ][9]<=-127; ws[7][2 ][10]<= -46; ws[7][2 ][11]<=  74; ws[7][2 ][12]<= 151; ws[7][2 ][13]<= -43; ws[7][2 ][14]<=  68; ws[7][2 ][15]<= 219;
        ws[7][3 ][0]<= -41; ws[7][3 ][1]<= -90; ws[7][3 ][2]<= 120; ws[7][3 ][3]<=-338; ws[7][3 ][4]<=-459; ws[7][3 ][5]<=-181; ws[7][3 ][6]<=-163; ws[7][3 ][7]<= -87; ws[7][3 ][8]<=  86; ws[7][3 ][9]<=-147; ws[7][3 ][10]<= 155; ws[7][3 ][11]<=-228; ws[7][3 ][12]<=-204; ws[7][3 ][13]<=-129; ws[7][3 ][14]<= -19; ws[7][3 ][15]<= -87;
        ws[7][4 ][0]<= 145; ws[7][4 ][1]<= 133; ws[7][4 ][2]<= 225; ws[7][4 ][3]<= 151; ws[7][4 ][4]<=  21; ws[7][4 ][5]<=  66; ws[7][4 ][6]<= 116; ws[7][4 ][7]<=  52; ws[7][4 ][8]<=  88; ws[7][4 ][9]<=  69; ws[7][4 ][10]<= -51; ws[7][4 ][11]<= 168; ws[7][4 ][12]<= 201; ws[7][4 ][13]<=-217; ws[7][4 ][14]<= 109; ws[7][4 ][15]<= 131;
        ws[7][5 ][0]<= 380; ws[7][5 ][1]<= -54; ws[7][5 ][2]<=-163; ws[7][5 ][3]<= -85; ws[7][5 ][4]<=  36; ws[7][5 ][5]<=-207; ws[7][5 ][6]<=-203; ws[7][5 ][7]<= 149; ws[7][5 ][8]<=  -3; ws[7][5 ][9]<= -52; ws[7][5 ][10]<= -76; ws[7][5 ][11]<=-164; ws[7][5 ][12]<=-245; ws[7][5 ][13]<= 383; ws[7][5 ][14]<= 268; ws[7][5 ][15]<=-230;
        ws[7][6 ][0]<=-164; ws[7][6 ][1]<= -81; ws[7][6 ][2]<= -38; ws[7][6 ][3]<=  43; ws[7][6 ][4]<= 191; ws[7][6 ][5]<=  43; ws[7][6 ][6]<= -50; ws[7][6 ][7]<= 160; ws[7][6 ][8]<=-216; ws[7][6 ][9]<= -27; ws[7][6 ][10]<= 163; ws[7][6 ][11]<=  72; ws[7][6 ][12]<= -26; ws[7][6 ][13]<= 245; ws[7][6 ][14]<=-141; ws[7][6 ][15]<= -89;
        ws[7][7 ][0]<=  70; ws[7][7 ][1]<=-164; ws[7][7 ][2]<=-174; ws[7][7 ][3]<=-221; ws[7][7 ][4]<=   4; ws[7][7 ][5]<=-104; ws[7][7 ][6]<=-266; ws[7][7 ][7]<=  56; ws[7][7 ][8]<= 234; ws[7][7 ][9]<=-144; ws[7][7 ][10]<= 229; ws[7][7 ][11]<=-193; ws[7][7 ][12]<= -56; ws[7][7 ][13]<= -67; ws[7][7 ][14]<=  66; ws[7][7 ][15]<= -81;
        ws[7][8 ][0]<=   8; ws[7][8 ][1]<= 220; ws[7][8 ][2]<=-188; ws[7][8 ][3]<=  98; ws[7][8 ][4]<= 252; ws[7][8 ][5]<= 202; ws[7][8 ][6]<=  44; ws[7][8 ][7]<=  16; ws[7][8 ][8]<=  -7; ws[7][8 ][9]<= 288; ws[7][8 ][10]<=  31; ws[7][8 ][11]<=  62; ws[7][8 ][12]<=  15; ws[7][8 ][13]<= 193; ws[7][8 ][14]<=   2; ws[7][8 ][15]<= -47;
        ws[7][9 ][0]<= 199; ws[7][9 ][1]<= 181; ws[7][9 ][2]<=-133; ws[7][9 ][3]<=  40; ws[7][9 ][4]<= -38; ws[7][9 ][5]<= -23; ws[7][9 ][6]<=  47; ws[7][9 ][7]<=-182; ws[7][9 ][8]<= 326; ws[7][9 ][9]<= 159; ws[7][9 ][10]<=-277; ws[7][9 ][11]<= 143; ws[7][9 ][12]<= 147; ws[7][9 ][13]<=-249; ws[7][9 ][14]<= 171; ws[7][9 ][15]<=  76;
        ws[7][10][0]<= 130; ws[7][10][1]<=-196; ws[7][10][2]<= 174; ws[7][10][3]<= -29; ws[7][10][4]<=-106; ws[7][10][5]<=-110; ws[7][10][6]<= -98; ws[7][10][7]<= 184; ws[7][10][8]<=  29; ws[7][10][9]<=-233; ws[7][10][10]<= 158; ws[7][10][11]<=-176; ws[7][10][12]<=-154; ws[7][10][13]<= 241; ws[7][10][14]<= 127; ws[7][10][15]<=-172;
        ws[7][11][0]<=-103; ws[7][11][1]<= 275; ws[7][11][2]<= 156; ws[7][11][3]<= 233; ws[7][11][4]<=  17; ws[7][11][5]<=  12; ws[7][11][6]<= 272; ws[7][11][7]<=-275; ws[7][11][8]<= 142; ws[7][11][9]<= 213; ws[7][11][10]<=-174; ws[7][11][11]<= -55; ws[7][11][12]<= 124; ws[7][11][13]<= 128; ws[7][11][14]<= -32; ws[7][11][15]<= 212;
        ws[7][12][0]<= -94; ws[7][12][1]<= 157; ws[7][12][2]<= 147; ws[7][12][3]<= 189; ws[7][12][4]<=  69; ws[7][12][5]<= 108; ws[7][12][6]<= 130; ws[7][12][7]<=-456; ws[7][12][8]<=  95; ws[7][12][9]<= 103; ws[7][12][10]<=-175; ws[7][12][11]<= 250; ws[7][12][12]<= 290; ws[7][12][13]<=  35; ws[7][12][14]<=  33; ws[7][12][15]<= 154;
        ws[7][13][0]<= 245; ws[7][13][1]<= -19; ws[7][13][2]<= -34; ws[7][13][3]<= 209; ws[7][13][4]<=-114; ws[7][13][5]<=-233; ws[7][13][6]<=  88; ws[7][13][7]<=-211; ws[7][13][8]<= 390; ws[7][13][9]<= -87; ws[7][13][10]<=-226; ws[7][13][11]<= 131; ws[7][13][12]<= 227; ws[7][13][13]<= -84; ws[7][13][14]<= 250; ws[7][13][15]<=  41;
        ws[7][14][0]<= 277; ws[7][14][1]<=-162; ws[7][14][2]<=  13; ws[7][14][3]<=  40; ws[7][14][4]<= -61; ws[7][14][5]<=-157; ws[7][14][6]<=  13; ws[7][14][7]<= -53; ws[7][14][8]<=  60; ws[7][14][9]<=-224; ws[7][14][10]<= 232; ws[7][14][11]<=-141; ws[7][14][12]<=-153; ws[7][14][13]<= 469; ws[7][14][14]<= 215; ws[7][14][15]<= -56;
        ws[7][15][0]<= -80; ws[7][15][1]<=   1; ws[7][15][2]<= 401; ws[7][15][3]<= 117; ws[7][15][4]<=-135; ws[7][15][5]<= -42; ws[7][15][6]<= -58; ws[7][15][7]<=   5; ws[7][15][8]<= 323; ws[7][15][9]<=-233; ws[7][15][10]<=  77; ws[7][15][11]<= 142; ws[7][15][12]<= 296; ws[7][15][13]<= -17; ws[7][15][14]<= 339; ws[7][15][15]<= 172;
    end

    always@(posedge clk) begin
        if(rst) begin
            w    <=0;
            ready<=0;
        end else if(start) begin
            w    <=ws[layer_sel][input_filter][output_filter];
            ready<=1; 
        end
    end
endmodule