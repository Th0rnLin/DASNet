`timescale 1ns/ 1ps

module conv_encoder_weights_memory(
    input wire                clk,
    input wire                rst,
    input wire                start,
    input wire        [3: 0]  input_filter,  // 14
    input wire        [3: 0]  output_filter, // 16
    output reg signed [17: 0] w,
    output reg                ready
);
    reg signed [17: 0] ws [0: 13][0: 15];

    initial begin
        ws[0 ][0 ]<=  267; ws[0 ][1 ]<=  -20; ws[0 ][2 ]<=  151; ws[0 ][3 ]<=   35; ws[0 ][4 ]<= -141;
        ws[0 ][5 ]<=   48; ws[0 ][6 ]<=  408; ws[0 ][7 ]<= -172; ws[0 ][8 ]<=  -80; ws[0 ][9 ]<=  151;
        ws[0 ][10]<=   87; ws[0 ][11]<= -169; ws[0 ][12]<=   58; ws[0 ][13]<= -103; ws[0 ][14]<=  156;
        ws[0 ][15]<= -148;
        ws[1 ][0 ]<=  -93; ws[1 ][1 ]<= -361; ws[1 ][2 ]<= -163; ws[1 ][3 ]<=   67; ws[1 ][4 ]<=  -51;
        ws[1 ][5 ]<= -192; ws[1 ][6 ]<=  229; ws[1 ][7 ]<=  237; ws[1 ][8 ]<=   33; ws[1 ][9 ]<= -301;
        ws[1 ][10]<= -340; ws[1 ][11]<=  -55; ws[1 ][12]<=  -48; ws[1 ][13]<= -288; ws[1 ][14]<=  305;
        ws[1 ][15]<=  240;
        ws[2 ][0 ]<=  -60; ws[2 ][1 ]<=  296; ws[2 ][2 ]<=-1570; ws[2 ][3 ]<=  701; ws[2 ][4 ]<=   10;
        ws[2 ][5 ]<=  698; ws[2 ][6 ]<=  855; ws[2 ][7 ]<=  880; ws[2 ][8 ]<= -886; ws[2 ][9 ]<=  389;
        ws[2 ][10]<=  862; ws[2 ][11]<= -129; ws[2 ][12]<=-1738; ws[2 ][13]<= -199; ws[2 ][14]<=-1090;
        ws[2 ][15]<= -921;
        ws[3 ][0 ]<=   39; ws[3 ][1 ]<= -108; ws[3 ][2 ]<=  285; ws[3 ][3 ]<= -190; ws[3 ][4 ]<= -112;
        ws[3 ][5 ]<=  -27; ws[3 ][6 ]<=  212; ws[3 ][7 ]<= -168; ws[3 ][8 ]<=  153; ws[3 ][9 ]<= -188;
        ws[3 ][10]<=  -40; ws[3 ][11]<=  -55; ws[3 ][12]<=   66; ws[3 ][13]<=  -44; ws[3 ][14]<=   51;
        ws[3 ][15]<= -110;
        ws[4 ][0 ]<=  139; ws[4 ][1 ]<= -182; ws[4 ][2 ]<=  -24; ws[4 ][3 ]<=  122; ws[4 ][4 ]<=  187;
        ws[4 ][5 ]<=  -70; ws[4 ][6 ]<=   66; ws[4 ][7 ]<=  172; ws[4 ][8 ]<=   13; ws[4 ][9 ]<=  -41;
        ws[4 ][10]<=   11; ws[4 ][11]<=  162; ws[4 ][12]<=   64; ws[4 ][13]<=  -18; ws[4 ][14]<=  -95;
        ws[4 ][15]<=  -90;
        ws[5 ][0 ]<=   46; ws[5 ][1 ]<=  119; ws[5 ][2 ]<=  -61; ws[5 ][3 ]<= -180; ws[5 ][4 ]<=  154;
        ws[5 ][5 ]<=  -29; ws[5 ][6 ]<=   44; ws[5 ][7 ]<= -162; ws[5 ][8 ]<=  171; ws[5 ][9 ]<= -127;
        ws[5 ][10]<=  -69; ws[5 ][11]<=   50; ws[5 ][12]<= -104; ws[5 ][13]<= -117; ws[5 ][14]<=  231;
        ws[5 ][15]<=  237;
        ws[6 ][0 ]<= -502; ws[6 ][1 ]<= -151; ws[6 ][2 ]<=  -39; ws[6 ][3 ]<=  523; ws[6 ][4 ]<= -603;
        ws[6 ][5 ]<=  678; ws[6 ][6 ]<=  490; ws[6 ][7 ]<= -189; ws[6 ][8 ]<=-1093; ws[6 ][9 ]<=  173;
        ws[6 ][10]<=  -47; ws[6 ][11]<= -766; ws[6 ][12]<=  -12; ws[6 ][13]<=  620; ws[6 ][14]<=  233;
        ws[6 ][15]<= -267;
        ws[7 ][0 ]<=  -94; ws[7 ][1 ]<=  -86; ws[7 ][2 ]<=  -70; ws[7 ][3 ]<=  -97; ws[7 ][4 ]<=   16;
        ws[7 ][5 ]<=   73; ws[7 ][6 ]<=  463; ws[7 ][7 ]<=  277; ws[7 ][8 ]<= -115; ws[7 ][9 ]<= -215;
        ws[7 ][10]<=   57; ws[7 ][11]<=  108; ws[7 ][12]<=  -89; ws[7 ][13]<= -158; ws[7 ][14]<= -158;
        ws[7 ][15]<=  178;
        ws[8 ][0 ]<=  303; ws[8 ][1 ]<= -199; ws[8 ][2 ]<=  120; ws[8 ][3 ]<=   78; ws[8 ][4 ]<= -181;
        ws[8 ][5 ]<=  -14; ws[8 ][6 ]<= -171; ws[8 ][7 ]<=   73; ws[8 ][8 ]<=   34; ws[8 ][9 ]<=  -33;
        ws[8 ][10]<=  327; ws[8 ][11]<=  309; ws[8 ][12]<=   66; ws[8 ][13]<= -107; ws[8 ][14]<=  -83;
        ws[8 ][15]<=    5;
        ws[9 ][0 ]<=  190; ws[9 ][1 ]<=  503; ws[9 ][2 ]<=  -58; ws[9 ][3 ]<=   62; ws[9 ][4 ]<=  393;
        ws[9 ][5 ]<=  418; ws[9 ][6 ]<=  819; ws[9 ][7 ]<=  450; ws[9 ][8 ]<= -859; ws[9 ][9 ]<= -153;
        ws[9 ][10]<=  585; ws[9 ][11]<=   90; ws[9 ][12]<= -460; ws[9 ][13]<=    2; ws[9 ][14]<= -568;
        ws[9 ][15]<= -899;
        ws[10][0 ]<= -290; ws[10][1 ]<=   15; ws[10][2 ]<=  112; ws[10][3 ]<=  -74; ws[10][4 ]<=  118;
        ws[10][5 ]<=  -89; ws[10][6 ]<=  108; ws[10][7 ]<=  -23; ws[10][8 ]<=   73; ws[10][9 ]<= -156;
        ws[10][10]<= -166; ws[10][11]<= -266; ws[10][12]<=   48; ws[10][13]<= -137; ws[10][14]<= -165;
        ws[10][15]<=  127;
        ws[11][0 ]<= -163; ws[11][1 ]<= -177; ws[11][2 ]<=   15; ws[11][3 ]<= -143; ws[11][4 ]<=  -46;
        ws[11][5 ]<=  101; ws[11][6 ]<= -100; ws[11][7 ]<= -196; ws[11][8 ]<=   -9; ws[11][9 ]<=   67;
        ws[11][10]<=  -31; ws[11][11]<=   92; ws[11][12]<=  -63; ws[11][13]<=  109; ws[11][14]<=   -6;
        ws[11][15]<=   62;
        ws[12][0 ]<= -110; ws[12][1 ]<= -156; ws[12][2 ]<=    1; ws[12][3 ]<=  -15; ws[12][4 ]<=  120;
        ws[12][5 ]<=   52; ws[12][6 ]<= -176; ws[12][7 ]<=  105; ws[12][8 ]<=   38; ws[12][9 ]<= -170;
        ws[12][10]<=   58; ws[12][11]<=  -11; ws[12][12]<=   51; ws[12][13]<= -251; ws[12][14]<=   50;
        ws[12][15]<=  374;
        ws[13][0 ]<= -373; ws[13][1 ]<= -586; ws[13][2 ]<=  156; ws[13][3 ]<=  390; ws[13][4 ]<= -432;
        ws[13][5 ]<=  518; ws[13][6 ]<= -147; ws[13][7 ]<= -165; ws[13][8 ]<= -934; ws[13][9 ]<=  352;
        ws[13][10]<= -180; ws[13][11]<=-1063; ws[13][12]<=   16; ws[13][13]<=  631; ws[13][14]<=  179;
        ws[13][15]<= -535;
    end

    always@(posedge clk) begin
        if(rst) begin
            w    <=0;
            ready<=0;
        end else if(start) begin
            w    <=ws[input_filter][output_filter];
            ready<=1; 
        end
    end
endmodule